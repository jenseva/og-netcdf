netcdf file:/Users/sevadjian/projects/og-netcdf/nc_out_2022_11_21.nc {
  dimensions:
    N_MEASUREMENTS = 24917;
    trajectory = 1;
  variables:
    int trajectory(trajectory=1);
      :cf_role = "trajectory_id";

    double TIME(N_MEASUREMENTS=24917);
      :axis = "T";
      :units = "seconds since 1970-01-01 00:00:00 UTC";
      :calendar = "julian";
      :standard_name = "time";
      :_fillValue = "-9999.0";
      :long_name = "Time";

    double LATITUDE(N_MEASUREMENTS=24917);
      :long_name = "Latitude";
      :standard_name = "latitude";
      :axis = "Y";
      :units = "degrees_north";

    double LONGITUDE(N_MEASUREMENTS=24917);
      :standard_name = "longitude";
      :axis = "X";
      :units = "degrees_east";
      :long_name = "Longitude";

    float DEPTH(N_MEASUREMENTS=24917);
      :units = "m";
      :positive = "Down";
      :axis = "Z";
      :long_name = "Depth";
      :standard_name = "Depth";

    double CHLA(N_MEASUREMENTS=24917);
      :_FillValue = NaN; // double
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water";
      :long_name = "Chlorophyll-a concentration";
      :units = "mg/m3";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :ancillary_variables = "CHLA_INSTRUMENT";

    float DENSITY(N_MEASUREMENTS=24917);
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :long_name = "Sea Water Density";
      :units = "kg m-3";
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :standard_name = "sea_water_density";
      :_FillValue = NaNf; // float

    double DOXY(N_MEASUREMENTS=24917);
      :_FillValue = NaN; // double
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water";
      :long_name = "Dissolved oxygen";
      :units = "micromol kg-1";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :ancillary_variables = "DOXY_QC DOXY_INSTRUMENT";

    byte DOXY_QC(N_MEASUREMENTS=24917);
      :long_name = "dissolved_oxygen Quality Flag";
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";

    int CHLA_INSTRUMENT(trajectory=1);
      :vocabulary = "https://docs.google.com/document/d/1dN90xkw9oCbLs0sPPhOmszdOjLpwcqxiK5mjeZP7abA/edit";
      :make_model = "ECO_FL";

    int DOXY_INSTRUMENT(trajectory=1);
      :vocabulary = "https://docs.google.com/document/d/1dN90xkw9oCbLs0sPPhOmszdOjLpwcqxiK5mjeZP7abA/edit";
      :make_model = "SEABIRD_SBE43F_IDO";

  // global attributes:
  :acknowledgement = "Funded by National Oceanic and Atmospheric Administration (NOAA): Global Ocean Monitoring and Observing (GOMO) Program, and Integrated Ocean Observing System. Supported by Instrument Development Group - Scripps Institution of Oceanography";
  :contributor_name = "Daniel Rudnick, Guilherme Castelao";
  :contributor_role = "Principal Investigator, Data Curator";
  :Conventions = "Unidata Dataset Discovery v1.0, COARDS, CF-1.6";
  :creator_email = "idgdata@ucsd.edu";
  :creator_institution = "University of California - San Diego; Scripps Institution of Oceanography";
  :creator_name = "Instrument Development Group";
  :creator_type = "group";
  :creator_url = "http://spraydata.ucsd.edu";
  :ctd_make_model = "Sea-Bird 41CP";
  :date_created = "2022-11-21T16:20:33.657126";
  :date_issued = "2022-11-21T16:20:40.338955";
  :date_modified = "2022-11-21T16:20:35.145640";
  :doi = "10.21238/S8SPRAY1618";
  :Easternmost_Easting = -123.336075; // double
  :format_version = "IOOS_Glider_NetCDF_v3.0.nc";
  :geospatial_bounds = "POLYGON ((-124.8602 37.761, -124.8303 37.7693, -124.852725 37.763075, -124.8602 37.761))";
  :geospatial_bounds_crs = "EPSG:4326";
  :geospatial_bounds_vertical_crs = "EPSG:5831";
  :geospatial_lat_max = 38.499936; // double
  :geospatial_lat_min = 37.2479; // double
  :geospatial_lat_units = "degrees_north";
  :geospatial_lon_max = -123.336075; // double
  :geospatial_lon_min = -126.1781; // double
  :geospatial_lon_units = "degrees_east";
  :geospatial_vertical_max = 504.1569f; // float
  :geospatial_vertical_min = 0.5955232f; // float
  :geospatial_vertical_positive = "down";
  :geospatial_vertical_units = "m";
  :gts_ingest = "true";
  :history = "readsat - 2022-11-21T08:20:25Z, fixgps3 - 2022-11-21T08:20:25Z, calcvelsat - 2022-11-21T08:20:25Z, autoqcctd - 2022-11-21T08:20:25Z, calox - 2022-11-21T08:20:26Z, calfchl - 2022-11-21T08:20:28Z, adpsat - 2022-11-21T08:20:32Z\n2022-11-21T18:23:47Z (local files)\n2022-11-21T18:23:47Z https://gliders.ioos.us/erddap/tabledap/sp011-20221014T1612.ncCF";
  :id = "sp011-20221014T1612";
  :infoUrl = "https://gliders.ioos.us/erddap/";
  :institution = "Scripps Institution of Oceanography";
  :instrument = "Sea-Bird 41CP";
  :ioos_dac_checksum = "d41d8cd98f00b204e9800998ecf8427e";
  :ioos_dac_completed = "False";
  :keywords = "AUVS > Autonomous Underwater Vehicles, Earth Science > Oceans > Ocean Pressure > Water Pressure, Earth Science > Oceans > Ocean Temperature > Water Temperature, Earth Science > Oceans > Salinity/Density > Conductivity, Earth Science > Oceans > Salinity/Density > Density, Earth Science > Oceans > Salinity/Density > Salinity, glider, In Situ Ocean-based platforms > Seaglider, Slocum, Spray, trajectory, underwater glider, water, wmo";
  :keywords_vocabulary = "GCMD Science Keywords";
  :license = "Creative Commons Attribution 4.0 International Public License (https://creativecommons.org/licenses/by/4.0/)";
  :Metadata_Conventions = "Unidata Dataset Discovery v1.0, COARDS, CF-1.6";
  :metadata_link = "http://spraydata.ucsd.edu";
  :naming_authority = "edu.ucsd.scripps";
  :network = "California Underwater Glider Network";
  :Northernmost_Northing = 38.499936; // double
  :platform = "sp011";
  :platform_institution = "Scripps";
  :platform_type = "Spray Glider";
  :processing_level = "Automatic quality control procedures were applied. For maximum quality assurance, use the delayed mode version of this dataset once it is available.";
  :product_version = "v3";
  :project = "California Underwater Glider Network - Line 56";
  :publisher_email = "idgdata@ucsd.edu";
  :publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography";
  :publisher_name = "Instrument Development Group";
  :publisher_type = "group";
  :publisher_url = "https://spraydata.ucsd.edu";
  :references = "Rudnick, D. L. (2016). Ocean research enabled by underwater gliders. Annual review of marine science, 8, 519-541, doi:10.1146/annurev-marine-122414-033913\n Rudnick, D. L., Davis, R. E., & Sherman, J. T. (2016). Spray Underwater Glider Operations. Journal of Atmospheric and Oceanic Technology, 33(6), 1113-1122, doi:10.1175/JTECH-D-15-0252.1\n Rudnick, D. L., Davis, R. E., Eriksen, C. C., Fratantoni, D. M., & Perry, M. J. (2004). Underwater gliders for ocean research. Marine Technology Society Journal, 38(2), 73-84, doi:10.4031/002533204787522703\n Sherman, J., Davis, R. E., Owens, W. B., & Valdes, J. (2001). The autonomous underwater glider \'Spray\'. IEEE Journal of oceanic Engineering, 26(4), 437-446, doi:10.1109/48.972076";
  :sea_name = "Coastal Waters of California";
  :site = "CUGN line 56";
  :source = "Observational data from a profiling underwater glider.";
  :sourceUrl = "(local files)";
  :Southernmost_Northing = 37.2479; // double
  :standard_name_vocabulary = "CF Standard Name Table v75";
  :subsetVariables = "wmo_id,trajectory,profile_id,time,latitude,longitude";
  :summary = "The overarching goal of the California Underwater Glider Network is to sustain baseline observations of climate variability off the coast of California. The technical approach is to deploy autonomous underwater gliders in a network to provide real-time data.\nThe CUGN uses Spray underwater gliders making repeated dives from the surface to 500 m and back, repeating the cycle every 3 hours, and traveling 3 km in the horizontal during that time. The CUGN includes gliders on three of the traditional cross-shore CalCOFI lines: line 66.7 off Monterey Bay, line 80 off Point Conception, and line 90 off Dana Point.\n The glider missions typically last about 100 days, and cover over 2000 km, thus providing 4-6 sections on lines extending 300-500 km offshore. Since 2005 the CUGN has covered 200,000 km over ground in 28 glider-years, while doing 90,000 dives.";
  :time_coverage_end = "2022-11-21T09:59:15Z";
  :time_coverage_start = "2022-10-14T16:48:45Z";
  :title = "sp011-20221014T1612";
  :trajectory = "sp011-20221014T1612";
  :Westernmost_Easting = -126.1781; // double
  :xglider_type = "profileObs";
  :featureType = "trajectory";
  :cdm_data_type = "Trajectory";

  data:
    trajectory = 
      {1}
    TIME = 
      {1.665763921E9, 1.665765846E9, 1.665765853E9, 1.665765861E9, 1.665765869E9, 1.665765877E9, 1.665765885E9, 1.665765893E9, 1.665765901E9, 1.665765909E9, 1.665765917E9, 1.665765925E9, 1.665765933E9, 1.665765941E9, 1.665765949E9, 1.665765957E9, 1.665765965E9, 1.665765973E9, 1.665765981E9, 1.665765989E9, 1.665765997E9, 1.665766005E9, 1.665766013E9, 1.665766021E9, 1.665766029E9, 1.665766037E9, 1.665766045E9, 1.665766053E9, 1.665766061E9, 1.665766069E9, 1.665766077E9, 1.665766085E9, 1.665766093E9, 1.665766101E9, 1.665766109E9, 1.665766117E9, 1.665766125E9, 1.665766133E9, 1.665766141E9, 1.665766149E9, 1.665766157E9, 1.665766165E9, 1.665766173E9, 1.665766181E9, 1.665766189E9, 1.665766197E9, 1.665766205E9, 1.665766213E9, 1.665766221E9, 1.665766229E9, 1.665766237E9, 1.665766245E9, 1.665766253E9, 1.665766261E9, 1.665766269E9, 1.665766277E9, 1.665766285E9, 1.665766293E9, 1.665766301E9, 1.665766309E9, 1.665766317E9, 1.665766325E9, 1.665766333E9, 1.665766341E9, 1.665766349E9, 1.665766357E9, 1.665766365E9, 1.665766373E9, 1.665766381E9, 1.665766389E9, 1.665766397E9, 1.665766405E9, 1.665766413E9, 1.665766421E9, 1.665766429E9, 1.665766437E9, 1.665766445E9, 1.665766453E9, 1.665766461E9, 1.665766469E9, 1.66576686E9, 1.66576704E9, 1.665768869E9, 1.665768877E9, 1.665768885E9, 1.665768893E9, 1.665768901E9, 1.665768909E9, 1.665768917E9, 1.665768925E9, 1.665768933E9, 1.665768941E9, 1.665768949E9, 1.665768957E9, 1.665768965E9, 1.665768973E9, 1.665768981E9, 1.665768989E9, 1.665768997E9, 1.665769005E9, 1.665769013E9, 1.665769021E9, 1.665769029E9, 1.665769037E9, 1.665769045E9, 1.665769053E9, 1.665769061E9, 1.665769069E9, 1.665769077E9, 1.665769085E9, 1.665769093E9, 1.665769101E9, 1.665769109E9, 1.665769117E9, 1.665769125E9, 1.665769133E9, 1.665769141E9, 1.665769149E9, 1.665769157E9, 1.665769165E9, 1.665769173E9, 1.665769181E9, 1.665769189E9, 1.665769197E9, 1.665769205E9, 1.665769213E9, 1.665769221E9, 1.665769229E9, 1.665769237E9, 1.665769245E9, 1.665769253E9, 1.665769261E9, 1.665769269E9, 1.665769277E9, 1.665769285E9, 1.665769293E9, 1.665769301E9, 1.665769309E9, 1.665769317E9, 1.665769325E9, 1.665769333E9, 1.665769341E9, 1.665769349E9, 1.665769357E9, 1.665769365E9, 1.665769373E9, 1.665769381E9, 1.665769389E9, 1.665769397E9, 1.665769405E9, 1.665769413E9, 1.665769421E9, 1.665769429E9, 1.665769437E9, 1.665769445E9, 1.665769453E9, 1.665769461E9, 1.665769469E9, 1.665769477E9, 1.665769485E9, 1.665769493E9, 1.665769501E9, 1.665769509E9, 1.66576974E9, 1.66576992E9, 1.665771884E9, 1.6657719E9, 1.665771916E9, 1.665771932E9, 1.665771948E9, 1.665771964E9, 1.66577198E9, 1.665771996E9, 1.665772012E9, 1.665772028E9, 1.665772044E9, 1.66577206E9, 1.665772076E9, 1.665772092E9, 1.665772108E9, 1.665772124E9, 1.66577214E9, 1.665772156E9, 1.665772172E9, 1.665772188E9, 1.665772204E9, 1.66577222E9, 1.665772236E9, 1.665772252E9, 1.665772268E9, 1.665772284E9, 1.6657723E9, 1.665772316E9, 1.665772332E9, 1.665772348E9, 1.665772364E9, 1.66577238E9, 1.665772396E9, 1.665772412E9, 1.665772428E9, 1.665772444E9, 1.66577246E9, 1.665772476E9, 1.665772492E9, 1.665772508E9, 1.665772524E9, 1.66577254E9, 1.665772556E9, 1.665772572E9, 1.665772588E9, 1.665772604E9, 1.66577262E9, 1.66577286E9, 1.66577304E9, 1.665775015E9, 1.665775031E9, 1.665775047E9, 1.665775063E9, 1.665775079E9, 1.665775095E9, 1.665775111E9, 1.665775127E9, 1.665775143E9, 1.665775159E9, 1.665775175E9, 1.665775191E9, 1.665775207E9, 1.665775223E9, 1.665775239E9, 1.665775255E9, 1.665775271E9, 1.665775287E9, 1.665775303E9, 1.665775319E9, 1.665775335E9, 1.665775351E9, 1.665775367E9, 1.665775383E9, 1.665775399E9, 1.665775415E9, 1.665775431E9, 1.665775447E9, 1.665775463E9, 1.665775479E9, 1.665775495E9, 1.665775511E9, 1.665775527E9, 1.665775543E9, 1.665775559E9, 1.665775575E9, 1.665775591E9, 1.665775607E9, 1.665775623E9, 1.665775639E9, 1.665775655E9, 1.665775671E9, 1.665775687E9, 1.665775703E9, 1.665775719E9, 1.665775735E9, 1.665775751E9, 1.665775767E9, 1.665775783E9, 1.665775799E9, 1.66577604E9, 1.66577622E9, 1.665778284E9, 1.6657783E9, 1.665778316E9, 1.665778332E9, 1.665778348E9, 1.665778364E9, 1.66577838E9, 1.665778396E9, 1.665778412E9, 1.665778428E9, 1.665778444E9, 1.66577846E9, 1.665778476E9, 1.665778492E9, 1.665778508E9, 1.665778524E9, 1.66577854E9, 1.665778556E9, 1.665778572E9, 1.665778588E9, 1.665778604E9, 1.66577862E9, 1.665778636E9, 1.665778652E9, 1.665778668E9, 1.665778684E9, 1.6657787E9, 1.665778716E9, 1.665778732E9, 1.665778748E9, 1.665778764E9, 1.66577878E9, 1.665778796E9, 1.665778812E9, 1.665778828E9, 1.665778844E9, 1.66577886E9, 1.665778876E9, 1.665778892E9, 1.665778908E9, 1.665778924E9, 1.66577894E9, 1.665778956E9, 1.665778972E9, 1.665778988E9, 1.665779004E9, 1.66577902E9, 1.665779036E9, 1.665779052E9, 1.665779068E9, 1.665779084E9, 1.6657791E9, 1.66577934E9, 1.66577952E9, 1.66578158E9, 1.665781596E9, 1.665781612E9, 1.665781628E9, 1.665781644E9, 1.66578166E9, 1.665781676E9, 1.665781692E9, 1.665781708E9, 1.665781724E9, 1.66578174E9, 1.665781756E9, 1.665781772E9, 1.665781788E9, 1.665781804E9, 1.66578182E9, 1.665781836E9, 1.665781852E9, 1.665781868E9, 1.665781884E9, 1.6657819E9, 1.665781916E9, 1.665781932E9, 1.665781948E9, 1.665781964E9, 1.66578198E9, 1.665781996E9, 1.665782012E9, 1.665782028E9, 1.665782044E9, 1.66578206E9, 1.665782076E9, 1.665782092E9, 1.665782108E9, 1.665782124E9, 1.66578214E9, 1.665782156E9, 1.665782172E9, 1.665782188E9, 1.665782204E9, 1.66578222E9, 1.665782236E9, 1.665782252E9, 1.665782268E9, 1.665782284E9, 1.6657823E9, 1.665782316E9, 1.665782332E9, 1.665782348E9, 1.665782364E9, 1.66578238E9, 1.665782396E9, 1.665782412E9, 1.665782428E9, 1.665782444E9, 1.66578246E9, 1.6657827E9, 1.66578294E9, 1.665784999E9, 1.665785015E9, 1.665785031E9, 1.665785047E9, 1.665785063E9, 1.665785079E9, 1.665785095E9, 1.665785111E9, 1.665785127E9, 1.665785143E9, 1.665785159E9, 1.665785175E9, 1.665785191E9, 1.665785207E9, 1.665785223E9, 1.665785239E9, 1.665785255E9, 1.665785271E9, 1.665785287E9, 1.665785303E9, 1.665785319E9, 1.665785335E9, 1.665785351E9, 1.665785367E9, 1.665785383E9, 1.665785399E9, 1.665785415E9, 1.665785431E9, 1.665785447E9, 1.665785463E9, 1.665785479E9, 1.665785495E9, 1.665785511E9, 1.665785527E9, 1.665785543E9, 1.665785559E9, 1.665785575E9, 1.665785591E9, 1.665785607E9, 1.665785623E9, 1.665785639E9, 1.665785655E9, 1.665785671E9, 1.665785687E9, 1.665785703E9, 1.665785719E9, 1.665785735E9, 1.665785751E9, 1.665785767E9, 1.665785783E9, 1.665785799E9, 1.665785815E9, 1.665785831E9, 1.665785847E9, 1.665785863E9, 1.665785879E9, 1.66578612E9, 1.6657863E9, 1.665788419E9, 1.665788435E9, 1.665788451E9, 1.665788467E9, 1.665788483E9, 1.665788499E9, 1.665788515E9, 1.665788531E9, 1.665788547E9, 1.665788563E9, 1.665788579E9, 1.665788595E9, 1.665788611E9, 1.665788627E9, 1.665788643E9, 1.665788659E9, 1.665788675E9, 1.665788691E9, 1.665788707E9, 1.665788723E9, 1.665788739E9, 1.665788755E9, 1.665788771E9, 1.665788787E9, 1.665788803E9, 1.665788819E9, 1.665788835E9, 1.665788851E9, 1.665788867E9, 1.665788883E9, 1.665788899E9, 1.665788915E9, 1.665788931E9, 1.665788947E9, 1.665788963E9, 1.665788979E9, 1.665788995E9, 1.665789011E9, 1.665789027E9, 1.665789043E9, 1.665789059E9, 1.665789075E9, 1.665789091E9, 1.665789107E9, 1.665789123E9, 1.665789139E9, 1.665789155E9, 1.665789171E9, 1.665789187E9, 1.665789203E9, 1.665789219E9, 1.665789235E9, 1.665789251E9, 1.665789267E9, 1.665789283E9, 1.665789299E9, 1.66578954E9, 1.66578984E9, 1.665792025E9, 1.665792041E9, 1.665792057E9, 1.665792073E9, 1.665792089E9, 1.665792105E9, 1.665792121E9, 1.665792137E9, 1.665792153E9, 1.665792169E9, 1.665792185E9, 1.665792201E9, 1.665792217E9, 1.665792233E9, 1.665792249E9, 1.665792265E9, 1.665792281E9, 1.665792297E9, 1.665792313E9, 1.665792329E9, 1.665792345E9, 1.665792361E9, 1.665792377E9, 1.665792393E9, 1.665792409E9, 1.665792425E9, 1.665792441E9, 1.665792457E9, 1.665792473E9, 1.665792489E9, 1.665792505E9, 1.665792521E9, 1.665792537E9, 1.665792553E9, 1.665792569E9, 1.665792585E9, 1.665792601E9, 1.665792617E9, 1.665792633E9, 1.665792649E9, 1.665792665E9, 1.665792681E9, 1.665792697E9, 1.665792713E9, 1.665792729E9, 1.665792745E9, 1.665792761E9, 1.665792777E9, 1.665792793E9, 1.665792809E9, 1.665792825E9, 1.665792841E9, 1.665792857E9, 1.665792873E9, 1.665792889E9, 1.665792905E9, 1.665792921E9, 1.665792937E9, 1.665792953E9, 1.665792969E9, 1.6657932E9, 1.66579338E9, 1.665795583E9, 1.665795599E9, 1.665795615E9, 1.665795631E9, 1.665795647E9, 1.665795663E9, 1.665795679E9, 1.665795695E9, 1.665795711E9, 1.665795727E9, 1.665795743E9, 1.665795759E9, 1.665795775E9, 1.665795791E9, 1.665795807E9, 1.665795823E9, 1.665795839E9, 1.665795855E9, 1.665795871E9, 1.665795887E9, 1.665795903E9, 1.665795919E9, 1.665795935E9, 1.665795951E9, 1.665795967E9, 1.665795983E9, 1.665795999E9, 1.665796015E9, 1.665796031E9, 1.665796047E9, 1.665796063E9, 1.665796079E9, 1.665796095E9, 1.665796111E9, 1.665796127E9, 1.665796143E9, 1.665796159E9, 1.665796175E9, 1.665796191E9, 1.665796207E9, 1.665796223E9, 1.665796239E9, 1.665796255E9, 1.665796271E9, 1.665796287E9, 1.665796303E9, 1.665796319E9, 1.665796335E9, 1.665796351E9, 1.665796367E9, 1.665796383E9, 1.665796399E9, 1.665796415E9, 1.665796431E9, 1.665796447E9, 1.665796463E9, 1.665796479E9, 1.665796495E9, 1.665796511E9, 1.665796527E9, 1.665796543E9, 1.665796559E9, 1.6657968E9, 1.66579698E9, 1.665799364E9, 1.66579938E9, 1.665799396E9, 1.665799412E9, 1.665799428E9, 1.665799444E9, 1.66579946E9, 1.665799476E9, 1.665799492E9, 1.665799508E9, 1.665799524E9, 1.66579954E9, 1.665799556E9, 1.665799572E9, 1.665799588E9, 1.665799604E9, 1.66579962E9, 1.665799636E9, 1.665799652E9, 1.665799668E9, 1.665799684E9, 1.6657997E9, 1.665799716E9, 1.665799732E9, 1.665799748E9, 1.665799764E9, 1.66579978E9, 1.665799796E9, 1.665799812E9, 1.665799828E9, 1.665799844E9, 1.66579986E9, 1.665799876E9, 1.665799892E9, 1.665799908E9, 1.665799924E9, 1.66579994E9, 1.665799956E9, 1.665799972E9, 1.665799988E9, 1.665800004E9, 1.66580002E9, 1.665800036E9, 1.665800052E9, 1.665800068E9, 1.665800084E9, 1.6658001E9, 1.665800116E9, 1.665800132E9, 1.665800148E9, 1.665800164E9, 1.66580018E9, 1.665800196E9, 1.665800212E9, 1.665800228E9, 1.665800244E9, 1.66580026E9, 1.665800276E9, 1.665800292E9, 1.665800308E9, 1.665800324E9, 1.66580034E9, 1.66580058E9, 1.66580076E9, 1.6658032E9, 1.665803216E9, 1.665803232E9, 1.665803248E9, 1.665803264E9, 1.66580328E9, 1.665803296E9, 1.665803312E9, 1.665803328E9, 1.665803344E9, 1.66580336E9, 1.665803376E9, 1.665803392E9, 1.665803408E9, 1.665803424E9, 1.66580344E9, 1.665803456E9, 1.665803472E9, 1.665803488E9, 1.665803504E9, 1.66580352E9, 1.665803536E9, 1.665803552E9, 1.665803568E9, 1.665803584E9, 1.6658036E9, 1.665803616E9, 1.665803632E9, 1.665803648E9, 1.665803664E9, 1.66580368E9, 1.665803696E9, 1.665803712E9, 1.665803728E9, 1.665803744E9, 1.66580376E9, 1.665803776E9, 1.665803792E9, 1.665803808E9, 1.665803824E9, 1.66580384E9, 1.665803856E9, 1.665803872E9, 1.665803888E9, 1.665803904E9, 1.66580392E9, 1.665803936E9, 1.665803952E9, 1.665803968E9, 1.665803984E9, 1.665804E9, 1.665804016E9, 1.665804032E9, 1.665804048E9, 1.665804064E9, 1.66580408E9, 1.665804096E9, 1.665804112E9, 1.665804128E9, 1.665804144E9, 1.66580416E9, 1.665804176E9, 1.665804192E9, 1.665804208E9, 1.665804224E9, 1.66580424E9, 1.66580448E9, 1.66580466E9, 1.665807204E9, 1.665807236E9, 1.665807268E9, 1.6658073E9, 1.665807332E9, 1.665807364E9, 1.665807396E9, 1.665807428E9, 1.66580746E9, 1.665807492E9, 1.665807524E9, 1.665807556E9, 1.665807588E9, 1.66580762E9, 1.665807652E9, 1.665807684E9, 1.665807716E9, 1.665807748E9, 1.66580778E9, 1.665807812E9, 1.665807844E9, 1.665807876E9, 1.665807908E9, 1.66580794E9, 1.665807972E9, 1.665808004E9, 1.665808036E9, 1.665808068E9, 1.6658081E9, 1.665808132E9, 1.665808164E9, 1.665808196E9, 1.665808228E9, 1.66580826E9, 1.665808292E9, 1.665808324E9, 1.665808356E9, 1.665808388E9, 1.66580842E9, 1.66580868E9, 1.66580886E9, 1.665811562E9, 1.665811594E9, 1.665811626E9, 1.665811658E9, 1.66581169E9, 1.665811722E9, 1.665811754E9, 1.665811786E9, 1.665811818E9, 1.66581185E9, 1.665811882E9, 1.665811914E9, 1.665811946E9, 1.665811978E9, 1.66581201E9, 1.665812042E9, 1.665812074E9, 1.665812106E9, 1.665812138E9, 1.66581217E9, 1.665812202E9, 1.665812234E9, 1.665812266E9, 1.665812298E9, 1.66581233E9, 1.665812362E9, 1.665812394E9, 1.665812426E9, 1.665812458E9, 1.66581249E9, 1.665812522E9, 1.665812554E9, 1.665812586E9, 1.665812618E9, 1.66581265E9, 1.665812682E9, 1.665812714E9, 1.665812746E9, 1.665812778E9, 1.66581281E9, 1.66581306E9, 1.66581324E9, 1.665816252E9, 1.665816284E9, 1.665816316E9, 1.665816348E9, 1.66581638E9, 1.665816412E9, 1.665816444E9, 1.665816476E9, 1.665816508E9, 1.66581654E9, 1.665816572E9, 1.665816604E9, 1.665816636E9, 1.665816668E9, 1.6658167E9, 1.665816732E9, 1.665816764E9, 1.665816796E9, 1.665816828E9, 1.66581686E9, 1.665816892E9, 1.665816924E9, 1.665816956E9, 1.665816988E9, 1.66581702E9, 1.665817052E9, 1.665817084E9, 1.665817116E9, 1.665817148E9, 1.66581718E9, 1.665817212E9, 1.665817244E9, 1.665817276E9, 1.665817308E9, 1.66581734E9, 1.665817372E9, 1.665817404E9, 1.665817436E9, 1.665817468E9, 1.6658175E9, 1.665817532E9, 1.665817564E9, 1.665817596E9, 1.665817628E9, 1.66581766E9, 1.66581792E9, 1.6658181E9, 1.665821434E9, 1.665821466E9, 1.665821498E9, 1.66582153E9, 1.665821562E9, 1.665821594E9, 1.665821626E9, 1.665821658E9, 1.66582169E9, 1.665821722E9, 1.665821754E9, 1.665821786E9, 1.665821818E9, 1.66582185E9, 1.665821882E9, 1.665821914E9, 1.665821946E9, 1.665821978E9, 1.66582201E9, 1.665822042E9, 1.665822074E9, 1.665822106E9, 1.665822138E9, 1.66582217E9, 1.665822202E9, 1.665822234E9, 1.665822266E9, 1.665822298E9, 1.66582233E9, 1.665822362E9, 1.665822394E9, 1.665822426E9, 1.665822458E9, 1.66582249E9, 1.665822522E9, 1.665822554E9, 1.665822586E9, 1.665822618E9, 1.66582265E9, 1.665822682E9, 1.665822714E9, 1.665822746E9, 1.665822778E9, 1.66582281E9, 1.665822842E9, 1.665822874E9, 1.665822906E9, 1.665822938E9, 1.66582297E9, 1.665823002E9, 1.665823034E9, 1.665823066E9, 1.665823098E9, 1.66582313E9, 1.66582338E9, 1.66582356E9, 1.665827137E9, 1.665827169E9, 1.665827201E9, 1.665827233E9, 1.665827265E9, 1.665827297E9, 1.665827329E9, 1.665827361E9, 1.665827393E9, 1.665827425E9, 1.665827457E9, 1.665827489E9, 1.665827521E9, 1.665827553E9, 1.665827585E9, 1.665827617E9, 1.665827649E9, 1.665827681E9, 1.665827713E9, 1.665827745E9, 1.665827777E9, 1.665827809E9, 1.665827841E9, 1.665827873E9, 1.665827905E9, 1.665827937E9, 1.665827969E9, 1.665828001E9, 1.665828033E9, 1.665828065E9, 1.665828097E9, 1.665828129E9, 1.665828161E9, 1.665828193E9, 1.665828225E9, 1.665828257E9, 1.665828289E9, 1.665828321E9, 1.665828353E9, 1.665828385E9, 1.665828417E9, 1.665828449E9, 1.665828481E9, 1.665828513E9, 1.665828545E9, 1.665828577E9, 1.665828609E9, 1.665828641E9, 1.665828673E9, 1.665828705E9, 1.665828737E9, 1.665828769E9, 1.66582902E9, 1.6658292E9, 1.665832889E9, 1.665832921E9, 1.665832953E9, 1.665832985E9, 1.665833017E9, 1.665833049E9, 1.665833081E9, 1.665833113E9, 1.665833145E9, 1.665833177E9, 1.665833209E9, 1.665833241E9, 1.665833273E9, 1.665833305E9, 1.665833337E9, 1.665833369E9, 1.665833401E9, 1.665833433E9, 1.665833465E9, 1.665833497E9, 1.665833529E9, 1.665833561E9, 1.665833593E9, 1.665833625E9, 1.665833657E9, 1.665833689E9, 1.665833721E9, 1.665833753E9, 1.665833785E9, 1.665833817E9, 1.665833849E9, 1.665833881E9, 1.665833913E9, 1.665833945E9, 1.665833977E9, 1.665834009E9, 1.665834041E9, 1.665834073E9, 1.665834105E9, 1.665834137E9, 1.665834169E9, 1.665834201E9, 1.665834233E9, 1.665834265E9, 1.665834297E9, 1.665834329E9, 1.665834361E9, 1.665834393E9, 1.665834425E9, 1.665834457E9, 1.665834489E9, 1.665834521E9, 1.665834553E9, 1.665834585E9, 1.665834617E9, 1.665834649E9, 1.665834681E9, 1.665834713E9, 1.665834745E9, 1.665834777E9, 1.665834809E9, 1.66583508E9, 1.66583526E9, 1.66583941E9, 1.665839442E9, 1.665839474E9, 1.665839506E9, 1.665839538E9, 1.66583957E9, 1.665839602E9, 1.665839634E9, 1.665839666E9, 1.665839698E9, 1.66583973E9, 1.665839762E9, 1.665839794E9, 1.665839826E9, 1.665839858E9, 1.66583989E9, 1.665839922E9, 1.665839954E9, 1.665839986E9, 1.665840018E9, 1.66584005E9, 1.665840082E9, 1.665840114E9, 1.665840146E9, 1.665840178E9, 1.66584021E9, 1.665840242E9, 1.665840274E9, 1.665840306E9, 1.665840338E9, 1.66584037E9, 1.665840402E9, 1.665840434E9, 1.665840466E9, 1.665840498E9, 1.66584053E9, 1.665840562E9, 1.665840594E9, 1.665840626E9, 1.665840658E9, 1.66584069E9, 1.665840722E9, 1.665840754E9, 1.665840786E9, 1.665840818E9, 1.66584085E9, 1.665840882E9, 1.665840914E9, 1.665840946E9, 1.665840978E9, 1.66584101E9, 1.665841042E9, 1.665841074E9, 1.665841106E9, 1.665841138E9, 1.66584117E9, 1.665841202E9, 1.665841234E9, 1.665841266E9, 1.665841298E9, 1.66584133E9, 1.665841362E9, 1.665841394E9, 1.665841426E9, 1.665841458E9, 1.66584149E9, 1.665841522E9, 1.665841554E9, 1.665841586E9, 1.665841618E9, 1.66584165E9, 1.66584192E9, 1.6658421E9, 1.665846928E9, 1.66584696E9, 1.665846992E9, 1.665847024E9, 1.665847056E9, 1.665847088E9, 1.66584712E9, 1.665847152E9, 1.665847184E9, 1.665847216E9, 1.665847248E9, 1.66584728E9, 1.665847312E9, 1.665847344E9, 1.665847376E9, 1.665847408E9, 1.66584744E9, 1.665847472E9, 1.665847504E9, 1.665847536E9, 1.665847568E9, 1.6658476E9, 1.665847632E9, 1.665847664E9, 1.665847696E9, 1.665847728E9, 1.66584776E9, 1.665847792E9, 1.665847824E9, 1.665847856E9, 1.665847888E9, 1.66584792E9, 1.665847952E9, 1.665847984E9, 1.665848016E9, 1.665848048E9, 1.66584808E9, 1.665848112E9, 1.665848144E9, 1.665848176E9, 1.665848208E9, 1.66584824E9, 1.665848272E9, 1.665848304E9, 1.665848336E9, 1.665848368E9, 1.6658484E9, 1.665848432E9, 1.665848464E9, 1.665848496E9, 1.665848528E9, 1.66584856E9, 1.665848592E9, 1.665848624E9, 1.665848656E9, 1.665848688E9, 1.66584872E9, 1.665848752E9, 1.665848784E9, 1.665848816E9, 1.665848848E9, 1.66584888E9, 1.665848912E9, 1.665848944E9, 1.665848976E9, 1.665849008E9, 1.66584904E9, 1.665849072E9, 1.665849104E9, 1.665849136E9, 1.665849168E9, 1.6658492E9, 1.665849232E9, 1.665849264E9, 1.665849296E9, 1.665849328E9, 1.66584936E9, 1.66584966E9, 1.66584984E9, 1.66585462E9, 1.665854652E9, 1.665854684E9, 1.665854716E9, 1.665854748E9, 1.66585478E9, 1.665854812E9, 1.665854844E9, 1.665854876E9, 1.665854908E9, 1.66585494E9, 1.665854972E9, 1.665855004E9, 1.665855036E9, 1.665855068E9, 1.6658551E9, 1.665855132E9, 1.665855164E9, 1.665855196E9, 1.665855228E9, 1.66585526E9, 1.665855292E9, 1.665855324E9, 1.665855356E9, 1.665855388E9, 1.66585542E9, 1.665855452E9, 1.665855484E9, 1.665855516E9, 1.665855548E9, 1.66585558E9, 1.665855612E9, 1.665855644E9, 1.665855676E9, 1.665855708E9, 1.66585574E9, 1.665855772E9, 1.665855804E9, 1.665855836E9, 1.665855868E9, 1.6658559E9, 1.665855932E9, 1.665855964E9, 1.665855996E9, 1.665856028E9, 1.66585606E9, 1.665856092E9, 1.665856124E9, 1.665856156E9, 1.665856188E9, 1.66585622E9, 1.665856252E9, 1.665856284E9, 1.665856316E9, 1.665856348E9, 1.66585638E9, 1.665856412E9, 1.665856444E9, 1.665856476E9, 1.665856508E9, 1.66585654E9, 1.665856572E9, 1.665856604E9, 1.665856636E9, 1.665856668E9, 1.6658567E9, 1.665856732E9, 1.665856764E9, 1.665856796E9, 1.665856828E9, 1.66585686E9, 1.665856892E9, 1.665856924E9, 1.665856956E9, 1.665856988E9, 1.66585702E9, 1.665857052E9, 1.665857084E9, 1.665857116E9, 1.665857148E9, 1.66585718E9, 1.66585746E9, 1.66585776E9, 1.665862461E9, 1.665862493E9, 1.665862525E9, 1.665862557E9, 1.665862589E9, 1.665862621E9, 1.665862653E9, 1.665862685E9, 1.665862717E9, 1.665862749E9, 1.665862781E9, 1.665862813E9, 1.665862845E9, 1.665862877E9, 1.665862909E9, 1.665862941E9, 1.665862973E9, 1.665863005E9, 1.665863037E9, 1.665863069E9, 1.665863101E9, 1.665863133E9, 1.665863165E9, 1.665863197E9, 1.665863229E9, 1.665863261E9, 1.665863293E9, 1.665863325E9, 1.665863357E9, 1.665863389E9, 1.665863421E9, 1.665863453E9, 1.665863485E9, 1.665863517E9, 1.665863549E9, 1.665863581E9, 1.665863613E9, 1.665863645E9, 1.665863677E9, 1.665863709E9, 1.665863741E9, 1.665863773E9, 1.665863805E9, 1.665863837E9, 1.665863869E9, 1.665863901E9, 1.665863933E9, 1.665863965E9, 1.665863997E9, 1.665864029E9, 1.665864061E9, 1.665864093E9, 1.665864125E9, 1.665864157E9, 1.665864189E9, 1.665864221E9, 1.665864253E9, 1.665864285E9, 1.665864317E9, 1.665864349E9, 1.665864381E9, 1.665864413E9, 1.665864445E9, 1.665864477E9, 1.665864509E9, 1.665864541E9, 1.665864573E9, 1.665864605E9, 1.665864637E9, 1.665864669E9, 1.665864701E9, 1.665864733E9, 1.665864765E9, 1.665864797E9, 1.665864829E9, 1.665864861E9, 1.665864893E9, 1.665864925E9, 1.665864957E9, 1.665864989E9, 1.66586526E9, 1.66586544E9, 1.66587017E9, 1.665870202E9, 1.665870234E9, 1.665870266E9, 1.665870298E9, 1.66587033E9, 1.665870362E9, 1.665870394E9, 1.665870426E9, 1.665870458E9, 1.66587049E9, 1.665870522E9, 1.665870554E9, 1.665870586E9, 1.665870618E9, 1.66587065E9, 1.665870682E9, 1.665870714E9, 1.665870746E9, 1.665870778E9, 1.66587081E9, 1.665870842E9, 1.665870874E9, 1.665870906E9, 1.665870938E9, 1.66587097E9, 1.665871002E9, 1.665871034E9, 1.665871066E9, 1.665871098E9, 1.66587113E9, 1.665871162E9, 1.665871194E9, 1.665871226E9, 1.665871258E9, 1.66587129E9, 1.665871322E9, 1.665871354E9, 1.665871386E9, 1.665871418E9, 1.66587145E9, 1.665871482E9, 1.665871514E9, 1.665871546E9, 1.665871578E9, 1.66587161E9, 1.665871642E9, 1.665871674E9, 1.665871706E9, 1.665871738E9, 1.66587177E9, 1.665871802E9, 1.665871834E9, 1.665871866E9, 1.665871898E9, 1.66587193E9, 1.665871962E9, 1.665871994E9, 1.665872026E9, 1.665872058E9, 1.66587209E9, 1.665872122E9, 1.665872154E9, 1.665872186E9, 1.665872218E9, 1.66587225E9, 1.665872282E9, 1.665872314E9, 1.665872346E9, 1.665872378E9, 1.66587241E9, 1.665872442E9, 1.665872474E9, 1.665872506E9, 1.665872538E9, 1.66587257E9, 1.665872602E9, 1.665872634E9, 1.665872666E9, 1.665872698E9, 1.66587273E9, 1.665873E9, 1.66587318E9, 1.665878054E9, 1.665878086E9, 1.665878118E9, 1.66587815E9, 1.665878182E9, 1.665878214E9, 1.665878246E9, 1.665878278E9, 1.66587831E9, 1.665878342E9, 1.665878374E9, 1.665878406E9, 1.665878438E9, 1.66587847E9, 1.665878502E9, 1.665878534E9, 1.665878566E9, 1.665878598E9, 1.66587863E9, 1.665878662E9, 1.665878694E9, 1.665878726E9, 1.665878758E9, 1.66587879E9, 1.665878822E9, 1.665878854E9, 1.665878886E9, 1.665878918E9, 1.66587895E9, 1.665878982E9, 1.665879014E9, 1.665879046E9, 1.665879078E9, 1.66587911E9, 1.665879142E9, 1.665879174E9, 1.665879206E9, 1.665879238E9, 1.66587927E9, 1.665879302E9, 1.665879334E9, 1.665879366E9, 1.665879398E9, 1.66587943E9, 1.665879462E9, 1.665879494E9, 1.665879526E9, 1.665879558E9, 1.66587959E9, 1.665879622E9, 1.665879654E9, 1.665879686E9, 1.665879718E9, 1.66587975E9, 1.665879782E9, 1.665879814E9, 1.665879846E9, 1.665879878E9, 1.66587991E9, 1.665879942E9, 1.665879974E9, 1.665880006E9, 1.665880038E9, 1.66588007E9, 1.665880102E9, 1.665880134E9, 1.665880166E9, 1.665880198E9, 1.66588023E9, 1.665880262E9, 1.665880294E9, 1.665880326E9, 1.665880358E9, 1.66588039E9, 1.665880422E9, 1.665880454E9, 1.665880486E9, 1.665880518E9, 1.66588055E9, 1.665880582E9, 1.665880614E9, 1.665880646E9, 1.665880678E9, 1.66588071E9, 1.66588104E9, 1.66588128E9, 1.665886142E9, 1.665886174E9, 1.665886206E9, 1.665886238E9, 1.66588627E9, 1.665886302E9, 1.665886334E9, 1.665886366E9, 1.665886398E9, 1.66588643E9, 1.665886462E9, 1.665886494E9, 1.665886526E9, 1.665886558E9, 1.66588659E9, 1.665886622E9, 1.665886654E9, 1.665886686E9, 1.665886718E9, 1.66588675E9, 1.665886782E9, 1.665886814E9, 1.665886846E9, 1.665886878E9, 1.66588691E9, 1.665886942E9, 1.665886974E9, 1.665887006E9, 1.665887038E9, 1.66588707E9, 1.665887102E9, 1.665887134E9, 1.665887166E9, 1.665887198E9, 1.66588723E9, 1.665887262E9, 1.665887294E9, 1.665887326E9, 1.665887358E9, 1.66588739E9, 1.665887422E9, 1.665887454E9, 1.665887486E9, 1.665887518E9, 1.66588755E9, 1.665887582E9, 1.665887614E9, 1.665887646E9, 1.665887678E9, 1.66588771E9, 1.665887742E9, 1.665887774E9, 1.665887806E9, 1.665887838E9, 1.66588787E9, 1.665887902E9, 1.665887934E9, 1.665887966E9, 1.665887998E9, 1.66588803E9, 1.665888062E9, 1.665888094E9, 1.665888126E9, 1.665888158E9, 1.66588819E9, 1.665888222E9, 1.665888254E9, 1.665888286E9, 1.665888318E9, 1.66588835E9, 1.665888382E9, 1.665888414E9, 1.665888446E9, 1.665888478E9, 1.66588851E9, 1.665888542E9, 1.665888574E9, 1.665888606E9, 1.665888638E9, 1.66588867E9, 1.66588896E9, 1.66588914E9, 1.665894053E9, 1.665894085E9, 1.665894117E9, 1.665894149E9, 1.665894181E9, 1.665894213E9, 1.665894245E9, 1.665894277E9, 1.665894309E9, 1.665894341E9, 1.665894373E9, 1.665894405E9, 1.665894437E9, 1.665894469E9, 1.665894501E9, 1.665894533E9, 1.665894565E9, 1.665894597E9, 1.665894629E9, 1.665894661E9, 1.665894693E9, 1.665894725E9, 1.665894757E9, 1.665894789E9, 1.665894821E9, 1.665894853E9, 1.665894885E9, 1.665894917E9, 1.665894949E9, 1.665894981E9, 1.665895013E9, 1.665895045E9, 1.665895077E9, 1.665895109E9, 1.665895141E9, 1.665895173E9, 1.665895205E9, 1.665895237E9, 1.665895269E9, 1.665895301E9, 1.665895333E9, 1.665895365E9, 1.665895397E9, 1.665895429E9, 1.665895461E9, 1.665895493E9, 1.665895525E9, 1.665895557E9, 1.665895589E9, 1.665895621E9, 1.665895653E9, 1.665895685E9, 1.665895717E9, 1.665895749E9, 1.665895781E9, 1.665895813E9, 1.665895845E9, 1.665895877E9, 1.665895909E9, 1.665895941E9, 1.665895973E9, 1.665896005E9, 1.665896037E9, 1.665896069E9, 1.665896101E9, 1.665896133E9, 1.665896165E9, 1.665896197E9, 1.665896229E9, 1.665896261E9, 1.665896293E9, 1.665896325E9, 1.665896357E9, 1.665896389E9, 1.665896421E9, 1.665896453E9, 1.665896485E9, 1.665896517E9, 1.665896549E9, 1.665896581E9, 1.665896613E9, 1.665896645E9, 1.665896677E9, 1.665896709E9, 1.665896741E9, 1.665896773E9, 1.665896805E9, 1.665896837E9, 1.665896869E9, 1.66589718E9, 1.66589742E9, 1.665902236E9, 1.665902268E9, 1.6659023E9, 1.665902332E9, 1.665902364E9, 1.665902396E9, 1.665902428E9, 1.66590246E9, 1.665902492E9, 1.665902524E9, 1.665902556E9, 1.665902588E9, 1.66590262E9, 1.665902652E9, 1.665902684E9, 1.665902716E9, 1.665902748E9, 1.66590278E9, 1.665902812E9, 1.665902844E9, 1.665902876E9, 1.665902908E9, 1.66590294E9, 1.665902972E9, 1.665903004E9, 1.665903036E9, 1.665903068E9, 1.6659031E9, 1.665903132E9, 1.665903164E9, 1.665903196E9, 1.665903228E9, 1.66590326E9, 1.665903292E9, 1.665903324E9, 1.665903356E9, 1.665903388E9, 1.66590342E9, 1.665903452E9, 1.665903484E9, 1.665903516E9, 1.665903548E9, 1.66590358E9, 1.665903612E9, 1.665903644E9, 1.665903676E9, 1.665903708E9, 1.66590374E9, 1.665903772E9, 1.665903804E9, 1.665903836E9, 1.665903868E9, 1.6659039E9, 1.665903932E9, 1.665903964E9, 1.665903996E9, 1.665904028E9, 1.66590406E9, 1.665904092E9, 1.665904124E9, 1.665904156E9, 1.665904188E9, 1.66590422E9, 1.665904252E9, 1.665904284E9, 1.665904316E9, 1.665904348E9, 1.66590438E9, 1.665904412E9, 1.665904444E9, 1.665904476E9, 1.665904508E9, 1.66590454E9, 1.665904572E9, 1.665904604E9, 1.665904636E9, 1.665904668E9, 1.6659047E9, 1.665904732E9, 1.665904764E9, 1.665904796E9, 1.665904828E9, 1.66590486E9, 1.665904892E9, 1.665904924E9, 1.665904956E9, 1.665904988E9, 1.66590502E9, 1.66590534E9, 1.66590564E9, 1.66591048E9, 1.665910528E9, 1.665910576E9, 1.665910624E9, 1.665910672E9, 1.66591072E9, 1.665910768E9, 1.665910816E9, 1.665910864E9, 1.665910912E9, 1.66591096E9, 1.665911008E9, 1.665911056E9, 1.665911104E9, 1.665911152E9, 1.6659112E9, 1.665911248E9, 1.665911296E9, 1.665911344E9, 1.665911392E9, 1.66591144E9, 1.665911488E9, 1.665911536E9, 1.665911584E9, 1.665911632E9, 1.66591168E9, 1.665911728E9, 1.665911776E9, 1.665911824E9, 1.665911872E9, 1.66591192E9, 1.665911968E9, 1.665912016E9, 1.665912064E9, 1.665912112E9, 1.66591216E9, 1.665912208E9, 1.665912256E9, 1.665912304E9, 1.665912352E9, 1.6659124E9, 1.665912448E9, 1.665912496E9, 1.665912544E9, 1.665912592E9, 1.66591264E9, 1.665912688E9, 1.665912736E9, 1.665912784E9, 1.665912832E9, 1.66591288E9, 1.665912928E9, 1.665912976E9, 1.665913024E9, 1.665913072E9, 1.66591312E9, 1.665913168E9, 1.665913216E9, 1.665913264E9, 1.665913312E9, 1.66591336E9, 1.665913408E9, 1.665913456E9, 1.665913504E9, 1.665913552E9, 1.6659136E9, 1.665913648E9, 1.665913696E9, 1.665913744E9, 1.665913792E9, 1.66591384E9, 1.66591416E9, 1.66591434E9, 1.665917886E9, 1.665917934E9, 1.665917982E9, 1.66591803E9, 1.665918078E9, 1.665918126E9, 1.665918174E9, 1.665918222E9, 1.66591827E9, 1.665918318E9, 1.665918366E9, 1.665918414E9, 1.665918462E9, 1.66591851E9, 1.665918558E9, 1.665918606E9, 1.665918654E9, 1.665918702E9, 1.66591875E9, 1.665918798E9, 1.665918846E9, 1.665918894E9, 1.665918942E9, 1.66591899E9, 1.665919038E9, 1.665919086E9, 1.665919134E9, 1.665919182E9, 1.66591923E9, 1.665919278E9, 1.665919326E9, 1.665919374E9, 1.665919422E9, 1.66591947E9, 1.665919518E9, 1.665919566E9, 1.665919614E9, 1.665919662E9, 1.66591971E9, 1.665919758E9, 1.665919806E9, 1.665919854E9, 1.665919902E9, 1.66591995E9, 1.66592022E9, 1.6659204E9, 1.665923499E9, 1.665923547E9, 1.665923595E9, 1.665923643E9, 1.665923691E9, 1.665923739E9, 1.665923787E9, 1.665923835E9, 1.665923883E9, 1.665923931E9, 1.665923979E9, 1.665924027E9, 1.665924075E9, 1.665924123E9, 1.665924171E9, 1.665924219E9, 1.665924267E9, 1.665924315E9, 1.665924363E9, 1.665924411E9, 1.665924459E9, 1.665924507E9, 1.665924555E9, 1.665924603E9, 1.665924651E9, 1.665924699E9, 1.665924747E9, 1.665924795E9, 1.665924843E9, 1.665924891E9, 1.665924939E9, 1.6659252E9, 1.66592538E9, 1.665928043E9, 1.665928091E9, 1.665928139E9, 1.665928187E9, 1.665928235E9, 1.665928283E9, 1.665928331E9, 1.665928379E9, 1.665928427E9, 1.665928475E9, 1.665928523E9, 1.665928571E9, 1.665928619E9, 1.665928667E9, 1.665928715E9, 1.665928763E9, 1.665928811E9, 1.665928859E9, 1.665928907E9, 1.665928955E9, 1.665929003E9, 1.665929051E9, 1.665929099E9, 1.665929147E9, 1.665929195E9, 1.665929243E9, 1.665929291E9, 1.665929339E9, 1.66592958E9, 1.66592982E9, 1.665932448E9, 1.665932496E9, 1.665932544E9, 1.665932592E9, 1.66593264E9, 1.665932688E9, 1.665932736E9, 1.665932784E9, 1.665932832E9, 1.66593288E9, 1.665932928E9, 1.665932976E9, 1.665933024E9, 1.665933072E9, 1.66593312E9, 1.665933168E9, 1.665933216E9, 1.665933264E9, 1.665933312E9, 1.66593336E9, 1.665933408E9, 1.665933456E9, 1.665933504E9, 1.665933552E9, 1.6659336E9, 1.66593384E9, 1.66593402E9, 1.665936743E9, 1.665936791E9, 1.665936839E9, 1.665936887E9, 1.665936935E9, 1.665936983E9, 1.665937031E9, 1.665937079E9, 1.665937127E9, 1.665937175E9, 1.665937223E9, 1.665937271E9, 1.665937319E9, 1.665937367E9, 1.665937415E9, 1.665937463E9, 1.665937511E9, 1.665937559E9, 1.665937607E9, 1.665937655E9, 1.665937703E9, 1.665937751E9, 1.665937799E9, 1.66593804E9, 1.66593828E9, 1.665940847E9, 1.665940895E9, 1.665940943E9, 1.665940991E9, 1.665941039E9, 1.665941087E9, 1.665941135E9, 1.665941183E9, 1.665941231E9, 1.665941279E9, 1.665941327E9, 1.665941375E9, 1.665941423E9, 1.665941471E9, 1.665941519E9, 1.665941567E9, 1.665941615E9, 1.665941663E9, 1.665941711E9, 1.665941759E9, 1.665941807E9, 1.665941855E9, 1.665941903E9, 1.665941951E9, 1.665941999E9, 1.66594224E9, 1.66594248E9, 1.665945262E9, 1.66594531E9, 1.665945358E9, 1.665945406E9, 1.665945454E9, 1.665945502E9, 1.66594555E9, 1.665945598E9, 1.665945646E9, 1.665945694E9, 1.665945742E9, 1.66594579E9, 1.665945838E9, 1.665945886E9, 1.665945934E9, 1.665945982E9, 1.66594603E9, 1.665946078E9, 1.665946126E9, 1.665946174E9, 1.665946222E9, 1.66594627E9, 1.6659465E9, 1.66594674E9, 1.665948936E9, 1.665948984E9, 1.665949032E9, 1.66594908E9, 1.665949128E9, 1.665949176E9, 1.665949224E9, 1.665949272E9, 1.66594932E9, 1.665949368E9, 1.665949416E9, 1.665949464E9, 1.665949512E9, 1.66594956E9, 1.665949608E9, 1.665949656E9, 1.665949704E9, 1.665949752E9, 1.6659498E9, 1.665949848E9, 1.665949896E9, 1.665949944E9, 1.665949992E9, 1.66595004E9, 1.66595028E9, 1.66595046E9, 1.665952837E9, 1.665952885E9, 1.665952933E9, 1.665952981E9, 1.665953029E9, 1.665953077E9, 1.665953125E9, 1.665953173E9, 1.665953221E9, 1.665953269E9, 1.665953317E9, 1.665953365E9, 1.665953413E9, 1.665953461E9, 1.665953509E9, 1.665953557E9, 1.665953605E9, 1.665953653E9, 1.665953701E9, 1.665953749E9, 1.665953797E9, 1.665953845E9, 1.665953893E9, 1.665953941E9, 1.665953989E9, 1.66595424E9, 1.66595436E9, 1.665956676E9, 1.665956724E9, 1.665956772E9, 1.66595682E9, 1.665956868E9, 1.665956916E9, 1.665956964E9, 1.665957012E9, 1.66595706E9, 1.665957108E9, 1.665957156E9, 1.665957204E9, 1.665957252E9, 1.6659573E9, 1.665957348E9, 1.665957396E9, 1.665957444E9, 1.665957492E9, 1.66595754E9, 1.665957588E9, 1.665957636E9, 1.665957684E9, 1.665957732E9, 1.66595778E9, 1.66595802E9, 1.6659582E9, 1.665960564E9, 1.665960612E9, 1.66596066E9, 1.665960708E9, 1.665960756E9, 1.665960804E9, 1.665960852E9, 1.6659609E9, 1.665960948E9, 1.665960996E9, 1.665961044E9, 1.665961092E9, 1.66596114E9, 1.665961188E9, 1.665961236E9, 1.665961284E9, 1.665961332E9, 1.66596138E9, 1.665961428E9, 1.665961476E9, 1.665961524E9, 1.665961572E9, 1.66596162E9, 1.66596186E9, 1.66596216E9, 1.665964356E9, 1.665964404E9, 1.665964452E9, 1.6659645E9, 1.665964548E9, 1.665964596E9, 1.665964644E9, 1.665964692E9, 1.66596474E9, 1.665964788E9, 1.665964836E9, 1.665964884E9, 1.665964932E9, 1.66596498E9, 1.665965028E9, 1.665965076E9, 1.665965124E9, 1.665965172E9, 1.66596522E9, 1.66596546E9, 1.66596564E9, 1.665967682E9, 1.66596773E9, 1.665967778E9, 1.665967826E9, 1.665967874E9, 1.665967922E9, 1.66596797E9, 1.665968018E9, 1.665968066E9, 1.665968114E9, 1.665968162E9, 1.66596821E9, 1.665968258E9, 1.665968306E9, 1.665968354E9, 1.665968402E9, 1.66596845E9, 1.665968498E9, 1.665968546E9, 1.665968594E9, 1.665968642E9, 1.66596869E9, 1.66596894E9, 1.66596912E9, 1.665971179E9, 1.665971227E9, 1.665971275E9, 1.665971323E9, 1.665971371E9, 1.665971419E9, 1.665971467E9, 1.665971515E9, 1.665971563E9, 1.665971611E9, 1.665971659E9, 1.665971707E9, 1.665971755E9, 1.665971803E9, 1.665971851E9, 1.665971899E9, 1.66597212E9, 1.6659723E9, 1.665974252E9, 1.6659743E9, 1.665974348E9, 1.665974396E9, 1.665974444E9, 1.665974492E9, 1.66597454E9, 1.665974588E9, 1.665974636E9, 1.665974684E9, 1.665974732E9, 1.66597478E9, 1.665974828E9, 1.665974876E9, 1.665974924E9, 1.665974972E9, 1.66597502E9, 1.66597524E9, 1.66597542E9, 1.665977361E9, 1.665977409E9, 1.665977457E9, 1.665977505E9, 1.665977553E9, 1.665977601E9, 1.665977649E9, 1.665977697E9, 1.665977745E9, 1.665977793E9, 1.665977841E9, 1.665977889E9, 1.665977937E9, 1.665977985E9, 1.665978033E9, 1.665978081E9, 1.665978129E9, 1.66597836E9, 1.66597854E9, 1.665980424E9, 1.665980472E9, 1.66598052E9, 1.665980568E9, 1.665980616E9, 1.665980664E9, 1.665980712E9, 1.66598076E9, 1.665980808E9, 1.665980856E9, 1.665980904E9, 1.665980952E9, 1.665981E9, 1.665981048E9, 1.665981096E9, 1.665981144E9, 1.665981192E9, 1.66598124E9, 1.66598148E9, 1.66598166E9, 1.665983389E9, 1.665983437E9, 1.665983485E9, 1.665983533E9, 1.665983581E9, 1.665983629E9, 1.665983677E9, 1.665983725E9, 1.665983773E9, 1.665983821E9, 1.665983869E9, 1.665983917E9, 1.665983965E9, 1.665984013E9, 1.665984061E9, 1.665984109E9, 1.665984157E9, 1.665984205E9, 1.665984253E9, 1.665984301E9, 1.665984349E9, 1.6659846E9, 1.66598478E9, 1.665986577E9, 1.665986625E9, 1.665986673E9, 1.665986721E9, 1.665986769E9, 1.665986817E9, 1.665986865E9, 1.665986913E9, 1.665986961E9, 1.665987009E9, 1.665987057E9, 1.665987105E9, 1.665987153E9, 1.665987201E9, 1.665987249E9, 1.66598748E9, 1.66598766E9, 1.665989698E9, 1.665989746E9, 1.665989794E9, 1.665989842E9, 1.66598989E9, 1.665989938E9, 1.665989986E9, 1.665990034E9, 1.665990082E9, 1.66599013E9, 1.665990178E9, 1.665990226E9, 1.665990274E9, 1.665990322E9, 1.66599037E9, 1.6659906E9, 1.66599072E9, 1.665992997E9, 1.665993045E9, 1.665993093E9, 1.665993141E9, 1.665993189E9, 1.665993237E9, 1.665993285E9, 1.665993333E9, 1.665993381E9, 1.665993429E9, 1.665993477E9, 1.665993525E9, 1.665993573E9, 1.665993621E9, 1.665993669E9, 1.6659939E9, 1.66599408E9, 1.665995758E9, 1.665995806E9, 1.665995854E9, 1.665995902E9, 1.66599595E9, 1.665995998E9, 1.665996046E9, 1.665996094E9, 1.665996142E9, 1.66599619E9, 1.665996238E9, 1.665996286E9, 1.665996334E9, 1.665996382E9, 1.66599643E9, 1.66599666E9, 1.66599684E9, 1.66599853E9, 1.665998578E9, 1.665998626E9, 1.665998674E9, 1.665998722E9, 1.66599877E9, 1.665998818E9, 1.665998866E9, 1.665998914E9, 1.665998962E9, 1.66599901E9, 1.665999058E9, 1.665999106E9, 1.665999154E9, 1.665999202E9, 1.66599925E9, 1.66599948E9, 1.66599966E9, 1.666001841E9, 1.666001889E9, 1.666001937E9, 1.666001985E9, 1.666002033E9, 1.666002081E9, 1.666002129E9, 1.666002177E9, 1.666002225E9, 1.666002273E9, 1.666002321E9, 1.666002369E9, 1.666002417E9, 1.666002465E9, 1.666002513E9, 1.666002561E9, 1.666002609E9, 1.66600284E9, 1.66600302E9, 1.666004937E9, 1.666004985E9, 1.666005033E9, 1.666005081E9, 1.666005129E9, 1.666005177E9, 1.666005225E9, 1.666005273E9, 1.666005321E9, 1.666005369E9, 1.666005417E9, 1.666005465E9, 1.666005513E9, 1.666005561E9, 1.666005609E9, 1.66600584E9, 1.66600602E9, 1.66600784E9, 1.666007888E9, 1.666007936E9, 1.666007984E9, 1.666008032E9, 1.66600808E9, 1.666008128E9, 1.666008176E9, 1.666008224E9, 1.666008272E9, 1.66600832E9, 1.666008368E9, 1.666008416E9, 1.666008464E9, 1.666008512E9, 1.66600856E9, 1.66600878E9, 1.66600896E9, 1.666010626E9, 1.666010674E9, 1.666010722E9, 1.66601077E9, 1.666010818E9, 1.666010866E9, 1.666010914E9, 1.666010962E9, 1.66601101E9, 1.666011058E9, 1.666011106E9, 1.666011154E9, 1.666011202E9, 1.66601125E9, 1.66601148E9, 1.66601166E9, 1.666013565E9, 1.666013613E9, 1.666013661E9, 1.666013709E9, 1.666013757E9, 1.666013805E9, 1.666013853E9, 1.666013901E9, 1.666013949E9, 1.666013997E9, 1.666014045E9, 1.666014093E9, 1.666014141E9, 1.666014189E9, 1.66601442E9, 1.6660146E9, 1.666016529E9, 1.666016577E9, 1.666016625E9, 1.666016673E9, 1.666016721E9, 1.666016769E9, 1.666016817E9, 1.666016865E9, 1.666016913E9, 1.666016961E9, 1.666017009E9, 1.666017057E9, 1.666017105E9, 1.666017153E9, 1.666017201E9, 1.666017249E9, 1.66601748E9, 1.66601766E9, 1.666019446E9, 1.666019494E9, 1.666019542E9, 1.66601959E9, 1.666019638E9, 1.666019686E9, 1.666019734E9, 1.666019782E9, 1.66601983E9, 1.666019878E9, 1.666019926E9, 1.666019974E9, 1.666020022E9, 1.66602007E9, 1.6660203E9, 1.66602048E9, 1.666022266E9, 1.666022314E9, 1.666022362E9, 1.66602241E9, 1.666022458E9, 1.666022506E9, 1.666022554E9, 1.666022602E9, 1.66602265E9, 1.666022698E9, 1.666022746E9, 1.666022794E9, 1.666022842E9, 1.66602289E9, 1.66602312E9, 1.6660233E9, 1.666024976E9, 1.666025024E9, 1.666025072E9, 1.66602512E9, 1.666025168E9, 1.666025216E9, 1.666025264E9, 1.666025312E9, 1.66602536E9, 1.666025408E9, 1.666025456E9, 1.666025504E9, 1.666025552E9, 1.6660256E9, 1.66602582E9, 1.666026E9, 1.666027688E9, 1.666027736E9, 1.666027784E9, 1.666027832E9, 1.66602788E9, 1.666027928E9, 1.666027976E9, 1.666028024E9, 1.666028072E9, 1.66602812E9, 1.666028168E9, 1.666028216E9, 1.666028264E9, 1.666028312E9, 1.66602836E9, 1.66602858E9, 1.66602876E9, 1.666030556E9, 1.666030604E9, 1.666030652E9, 1.6660307E9, 1.666030748E9, 1.666030796E9, 1.666030844E9, 1.666030892E9, 1.66603094E9, 1.666030988E9, 1.666031036E9, 1.666031084E9, 1.666031132E9, 1.66603118E9, 1.6660314E9, 1.66603158E9, 1.666033178E9, 1.666033226E9, 1.666033274E9, 1.666033322E9, 1.66603337E9, 1.666033418E9, 1.666033466E9, 1.666033514E9, 1.666033562E9, 1.66603361E9, 1.666033658E9, 1.666033706E9, 1.666033754E9, 1.666033802E9, 1.66603385E9, 1.6660341E9, 1.66603428E9, 1.666035995E9, 1.666036043E9, 1.666036091E9, 1.666036139E9, 1.666036187E9, 1.666036235E9, 1.666036283E9, 1.666036331E9, 1.666036379E9, 1.666036427E9, 1.666036475E9, 1.666036523E9, 1.666036571E9, 1.666036619E9, 1.66603686E9, 1.6660371E9, 1.666037101E9, 1.666037102E9, 1.666037103E9, 1.666037104E9, 1.666037105E9, 1.666037106E9, 1.666037107E9, 1.666037108E9, 1.666037109E9, 1.66603711E9, 1.666037111E9, 1.666037112E9, 1.666037113E9, 1.666037114E9, 1.6660392E9, 1.666039201E9, 1.666040455E9, 1.666040503E9, 1.666040551E9, 1.666040599E9, 1.666040647E9, 1.666040695E9, 1.666040743E9, 1.666040791E9, 1.666040839E9, 1.666040887E9, 1.666040935E9, 1.666040983E9, 1.666041031E9, 1.666041079E9, 1.6660413E9, 1.66604148E9, 1.666041481E9, 1.666041482E9, 1.666041483E9, 1.666041484E9, 1.666041485E9, 1.666041486E9, 1.666041487E9, 1.666041488E9, 1.666041489E9, 1.66604149E9, 1.666041491E9, 1.666041492E9, 1.666041493E9, 1.666041494E9, 1.666041495E9, 1.666043747E9, 1.666043748E9, 1.666044812E9, 1.66604486E9, 1.666044908E9, 1.666044956E9, 1.666045004E9, 1.666045052E9, 1.6660451E9, 1.666045148E9, 1.666045196E9, 1.666045244E9, 1.666045292E9, 1.66604534E9, 1.66604556E9, 1.66604574E9, 1.666045741E9, 1.666045742E9, 1.666045743E9, 1.666045744E9, 1.666045745E9, 1.666045746E9, 1.666045747E9, 1.666045748E9, 1.666045749E9, 1.66604575E9, 1.666045751E9, 1.666045752E9, 1.666045753E9, 1.666045754E9, 1.666047905E9, 1.666047906E9, 1.666049011E9, 1.666049059E9, 1.666049107E9, 1.666049155E9, 1.666049203E9, 1.666049251E9, 1.666049299E9, 1.666049347E9, 1.666049395E9, 1.666049443E9, 1.666049491E9, 1.666049539E9, 1.66604976E9, 1.66604994E9, 1.666049941E9, 1.666049942E9, 1.666049943E9, 1.666049944E9, 1.666049945E9, 1.666049946E9, 1.666049947E9, 1.666049948E9, 1.666049949E9, 1.66604995E9, 1.666049951E9, 1.666049952E9, 1.666049953E9, 1.666049954E9, 1.666049955E9, 1.66605219E9, 1.666052191E9, 1.66605315E9, 1.666053198E9, 1.666053246E9, 1.666053294E9, 1.666053342E9, 1.66605339E9, 1.666053438E9, 1.666053486E9, 1.666053534E9, 1.666053582E9, 1.66605363E9, 1.66605384E9, 1.66605402E9, 1.666054021E9, 1.666054022E9, 1.666054023E9, 1.666054024E9, 1.666054025E9, 1.666054026E9, 1.666054027E9, 1.666054028E9, 1.666054029E9, 1.66605403E9, 1.666054031E9, 1.666054032E9, 1.666054033E9, 1.666054034E9, 1.666056271E9, 1.666056272E9, 1.66605732E9, 1.666057368E9, 1.666057416E9, 1.666057464E9, 1.666057512E9, 1.66605756E9, 1.666057608E9, 1.666057656E9, 1.666057704E9, 1.666057752E9, 1.6660578E9, 1.66605804E9, 1.66605822E9, 1.666058221E9, 1.666058222E9, 1.666058223E9, 1.666058224E9, 1.666058225E9, 1.666058226E9, 1.666058227E9, 1.666058228E9, 1.666058229E9, 1.66605823E9, 1.666058231E9, 1.666058232E9, 1.666058233E9, 1.66606023E9, 1.666060231E9, 1.666061433E9, 1.666061481E9, 1.666061529E9, 1.666061577E9, 1.666061625E9, 1.666061673E9, 1.666061721E9, 1.666061769E9, 1.666061817E9, 1.666061865E9, 1.666061913E9, 1.666061961E9, 1.666062009E9, 1.66606224E9, 1.66606248E9, 1.666062481E9, 1.666062482E9, 1.666062483E9, 1.666062484E9, 1.666062485E9, 1.666062486E9, 1.666062487E9, 1.666062488E9, 1.666062489E9, 1.66606249E9, 1.666062491E9, 1.666062492E9, 1.666062493E9, 1.666062494E9, 1.666064689E9, 1.66606469E9, 1.666065923E9, 1.666065971E9, 1.666066019E9, 1.666066067E9, 1.666066115E9, 1.666066163E9, 1.666066211E9, 1.666066259E9, 1.666066307E9, 1.666066355E9, 1.666066403E9, 1.666066451E9, 1.666066499E9, 1.66606674E9, 1.66606692E9, 1.666066921E9, 1.666066922E9, 1.666066923E9, 1.666066924E9, 1.666066925E9, 1.666066926E9, 1.666066927E9, 1.666066928E9, 1.666066929E9, 1.66606693E9, 1.666066931E9, 1.666066932E9, 1.666066933E9, 1.666066934E9, 1.666066935E9, 1.666069287E9, 1.666069288E9, 1.666070421E9, 1.666070469E9, 1.666070517E9, 1.666070565E9, 1.666070613E9, 1.666070661E9, 1.666070709E9, 1.666070757E9, 1.666070805E9, 1.666070853E9, 1.666070901E9, 1.666070949E9, 1.66607118E9, 1.66607142E9, 1.666073155E9, 1.666073203E9, 1.666073251E9, 1.666073299E9, 1.666073347E9, 1.666073395E9, 1.666073443E9, 1.666073491E9, 1.666073539E9, 1.666073587E9, 1.666073635E9, 1.666073683E9, 1.666073731E9, 1.666073779E9, 1.666074E9, 1.66607424E9, 1.666076018E9, 1.666076066E9, 1.666076114E9, 1.666076162E9, 1.66607621E9, 1.666076258E9, 1.666076306E9, 1.666076354E9, 1.666076402E9, 1.66607645E9, 1.666076498E9, 1.666076546E9, 1.666076594E9, 1.666076642E9, 1.66607669E9, 1.66607694E9, 1.66607712E9, 1.666078788E9, 1.666078836E9, 1.666078884E9, 1.666078932E9, 1.66607898E9, 1.666079028E9, 1.666079076E9, 1.666079124E9, 1.666079172E9, 1.66607922E9, 1.666079268E9, 1.666079316E9, 1.666079364E9, 1.666079412E9, 1.66607946E9, 1.6660797E9, 1.66607988E9, 1.666081676E9, 1.666081724E9, 1.666081772E9, 1.66608182E9, 1.666081868E9, 1.666081916E9, 1.666081964E9, 1.666082012E9, 1.66608206E9, 1.666082108E9, 1.666082156E9, 1.666082204E9, 1.666082252E9, 1.6660823E9, 1.66608252E9, 1.66608276E9, 1.666084485E9, 1.666084533E9, 1.666084581E9, 1.666084629E9, 1.666084677E9, 1.666084725E9, 1.666084773E9, 1.666084821E9, 1.666084869E9, 1.666084917E9, 1.666084965E9, 1.666085013E9, 1.666085061E9, 1.666085109E9, 1.66608534E9, 1.66608552E9, 1.666087317E9, 1.666087365E9, 1.666087413E9, 1.666087461E9, 1.666087509E9, 1.666087557E9, 1.666087605E9, 1.666087653E9, 1.666087701E9, 1.666087749E9, 1.666087797E9, 1.666087845E9, 1.666087893E9, 1.666087941E9, 1.666087989E9, 1.66608822E9, 1.6660884E9, 1.666090248E9, 1.666090296E9, 1.666090344E9, 1.666090392E9, 1.66609044E9, 1.666090488E9, 1.666090536E9, 1.666090584E9, 1.666090632E9, 1.66609068E9, 1.666090728E9, 1.666090776E9, 1.666090824E9, 1.666090872E9, 1.66609092E9, 1.66609116E9, 1.66609134E9, 1.666093281E9, 1.666093329E9, 1.666093377E9, 1.666093425E9, 1.666093473E9, 1.666093521E9, 1.666093569E9, 1.666093617E9, 1.666093665E9, 1.666093713E9, 1.666093761E9, 1.666093809E9, 1.666093857E9, 1.666093905E9, 1.666093953E9, 1.666094001E9, 1.666094049E9, 1.66609428E9, 1.66609458E9, 1.666096382E9, 1.66609643E9, 1.666096478E9, 1.666096526E9, 1.666096574E9, 1.666096622E9, 1.66609667E9, 1.666096718E9, 1.666096766E9, 1.666096814E9, 1.666096862E9, 1.66609691E9, 1.666096958E9, 1.666097006E9, 1.666097054E9, 1.666097102E9, 1.66609715E9, 1.6660974E9, 1.6660977E9, 1.66609963E9, 1.666099678E9, 1.666099726E9, 1.666099774E9, 1.666099822E9, 1.66609987E9, 1.666099918E9, 1.666099966E9, 1.666100014E9, 1.666100062E9, 1.66610011E9, 1.666100158E9, 1.666100206E9, 1.666100254E9, 1.666100302E9, 1.66610035E9, 1.66610058E9, 1.66610076E9, 1.6661027E9, 1.666102748E9, 1.666102796E9, 1.666102844E9, 1.666102892E9, 1.66610294E9, 1.666102988E9, 1.666103036E9, 1.666103084E9, 1.666103132E9, 1.66610318E9, 1.666103228E9, 1.666103276E9, 1.666103324E9, 1.666103372E9, 1.66610342E9, 1.66610364E9, 1.66610382E9, 1.66610575E9, 1.666105798E9, 1.666105846E9, 1.666105894E9, 1.666105942E9, 1.66610599E9, 1.666106038E9, 1.666106086E9, 1.666106134E9, 1.666106182E9, 1.66610623E9, 1.666106278E9, 1.666106326E9, 1.666106374E9, 1.666106422E9, 1.66610647E9, 1.6661067E9, 1.66610694E9, 1.666108931E9, 1.666108979E9, 1.666109027E9, 1.666109075E9, 1.666109123E9, 1.666109171E9, 1.666109219E9, 1.666109267E9, 1.666109315E9, 1.666109363E9, 1.666109411E9, 1.666109459E9, 1.666109507E9, 1.666109555E9, 1.666109603E9, 1.666109651E9, 1.666109699E9, 1.66610994E9, 1.66611018E9, 1.666112171E9, 1.666112219E9, 1.666112267E9, 1.666112315E9, 1.666112363E9, 1.666112411E9, 1.666112459E9, 1.666112507E9, 1.666112555E9, 1.666112603E9, 1.666112651E9, 1.666112699E9, 1.666112747E9, 1.666112795E9, 1.666112843E9, 1.666112891E9, 1.666112939E9, 1.66611318E9, 1.6661133E9, 1.666115292E9, 1.66611534E9, 1.666115388E9, 1.666115436E9, 1.666115484E9, 1.666115532E9, 1.66611558E9, 1.666115628E9, 1.666115676E9, 1.666115724E9, 1.666115772E9, 1.66611582E9, 1.666115868E9, 1.666115916E9, 1.666115964E9, 1.666116012E9, 1.66611606E9, 1.6661163E9, 1.66611648E9, 1.666118485E9, 1.666118533E9, 1.666118581E9, 1.666118629E9, 1.666118677E9, 1.666118725E9, 1.666118773E9, 1.666118821E9, 1.666118869E9, 1.666118917E9, 1.666118965E9, 1.666119013E9, 1.666119061E9, 1.666119109E9, 1.666119157E9, 1.666119205E9, 1.666119253E9, 1.666119301E9, 1.666119349E9, 1.6661196E9, 1.66611978E9, 1.666121845E9, 1.666121893E9, 1.666121941E9, 1.666121989E9, 1.666122037E9, 1.666122085E9, 1.666122133E9, 1.666122181E9, 1.666122229E9, 1.666122277E9, 1.666122325E9, 1.666122373E9, 1.666122421E9, 1.666122469E9, 1.666122517E9, 1.666122565E9, 1.666122613E9, 1.666122661E9, 1.666122709E9, 1.66612296E9, 1.66612314E9, 1.666125153E9, 1.666125201E9, 1.666125249E9, 1.666125297E9, 1.666125345E9, 1.666125393E9, 1.666125441E9, 1.666125489E9, 1.666125537E9, 1.666125585E9, 1.666125633E9, 1.666125681E9, 1.666125729E9, 1.666125777E9, 1.666125825E9, 1.666125873E9, 1.666125921E9, 1.666125969E9, 1.6661262E9, 1.66612644E9, 1.666128458E9, 1.666128506E9, 1.666128554E9, 1.666128602E9, 1.66612865E9, 1.666128698E9, 1.666128746E9, 1.666128794E9, 1.666128842E9, 1.66612889E9, 1.666128938E9, 1.666128986E9, 1.666129034E9, 1.666129082E9, 1.66612913E9, 1.666129178E9, 1.666129226E9, 1.666129274E9, 1.666129322E9, 1.66612937E9, 1.66612962E9, 1.6661298E9, 1.666131983E9, 1.666132031E9, 1.666132079E9, 1.666132127E9, 1.666132175E9, 1.666132223E9, 1.666132271E9, 1.666132319E9, 1.666132367E9, 1.666132415E9, 1.666132463E9, 1.666132511E9, 1.666132559E9, 1.666132607E9, 1.666132655E9, 1.666132703E9, 1.666132751E9, 1.666132799E9, 1.666132847E9, 1.666132895E9, 1.666132943E9, 1.666132991E9, 1.666133039E9, 1.66613328E9, 1.66613352E9, 1.666135761E9, 1.666135809E9, 1.666135857E9, 1.666135905E9, 1.666135953E9, 1.666136001E9, 1.666136049E9, 1.666136097E9, 1.666136145E9, 1.666136193E9, 1.666136241E9, 1.666136289E9, 1.666136337E9, 1.666136385E9, 1.666136433E9, 1.666136481E9, 1.666136529E9, 1.666136577E9, 1.666136625E9, 1.666136673E9, 1.666136721E9, 1.666136769E9, 1.666137E9, 1.66613718E9, 1.666139444E9, 1.666139492E9, 1.66613954E9, 1.666139588E9, 1.666139636E9, 1.666139684E9, 1.666139732E9, 1.66613978E9, 1.666139828E9, 1.666139876E9, 1.666139924E9, 1.666139972E9, 1.66614002E9, 1.666140068E9, 1.666140116E9, 1.666140164E9, 1.666140212E9, 1.66614026E9, 1.666140308E9, 1.666140356E9, 1.666140404E9, 1.666140452E9, 1.6661405E9, 1.66614078E9, 1.66614108E9, 1.666143475E9, 1.666143523E9, 1.666143571E9, 1.666143619E9, 1.666143667E9, 1.666143715E9, 1.666143763E9, 1.666143811E9, 1.666143859E9, 1.666143907E9, 1.666143955E9, 1.666144003E9, 1.666144051E9, 1.666144099E9, 1.666144147E9, 1.666144195E9, 1.666144243E9, 1.666144291E9, 1.666144339E9, 1.666144387E9, 1.666144435E9, 1.666144483E9, 1.666144531E9, 1.666144579E9, 1.66614486E9, 1.6661451E9, 1.666147478E9, 1.666147526E9, 1.666147574E9, 1.666147622E9, 1.66614767E9, 1.666147718E9, 1.666147766E9, 1.666147814E9, 1.666147862E9, 1.66614791E9, 1.666147958E9, 1.666148006E9, 1.666148054E9, 1.666148102E9, 1.66614815E9, 1.666148198E9, 1.666148246E9, 1.666148294E9, 1.666148342E9, 1.66614839E9, 1.666148438E9, 1.666148486E9, 1.666148534E9, 1.666148582E9, 1.66614863E9, 1.66614888E9, 1.66614906E9, 1.666151556E9, 1.666151604E9, 1.666151652E9, 1.6661517E9, 1.666151748E9, 1.666151796E9, 1.666151844E9, 1.666151892E9, 1.66615194E9, 1.666151988E9, 1.666152036E9, 1.666152084E9, 1.666152132E9, 1.66615218E9, 1.666152228E9, 1.666152276E9, 1.666152324E9, 1.666152372E9, 1.66615242E9, 1.666152468E9, 1.666152516E9, 1.666152564E9, 1.666152612E9, 1.66615266E9, 1.6661529E9, 1.66615308E9, 1.666155599E9, 1.666155647E9, 1.666155695E9, 1.666155743E9, 1.666155791E9, 1.666155839E9, 1.666155887E9, 1.666155935E9, 1.666155983E9, 1.666156031E9, 1.666156079E9, 1.666156127E9, 1.666156175E9, 1.666156223E9, 1.666156271E9, 1.666156319E9, 1.666156367E9, 1.666156415E9, 1.666156463E9, 1.666156511E9, 1.666156559E9, 1.666156607E9, 1.666156655E9, 1.666156703E9, 1.666156751E9, 1.666156799E9, 1.66615704E9, 1.66615722E9, 1.666159946E9, 1.666159994E9, 1.666160042E9, 1.66616009E9, 1.666160138E9, 1.666160186E9, 1.666160234E9, 1.666160282E9, 1.66616033E9, 1.666160378E9, 1.666160426E9, 1.666160474E9, 1.666160522E9, 1.66616057E9, 1.666160618E9, 1.666160666E9, 1.666160714E9, 1.666160762E9, 1.66616081E9, 1.666160858E9, 1.666160906E9, 1.666160954E9, 1.666161002E9, 1.66616105E9, 1.666161098E9, 1.666161146E9, 1.666161194E9, 1.666161242E9, 1.66616129E9, 1.66616154E9, 1.66616172E9, 1.666164681E9, 1.666164729E9, 1.666164777E9, 1.666164825E9, 1.666164873E9, 1.666164921E9, 1.666164969E9, 1.666165017E9, 1.666165065E9, 1.666165113E9, 1.666165161E9, 1.666165209E9, 1.666165257E9, 1.666165305E9, 1.666165353E9, 1.666165401E9, 1.666165449E9, 1.666165497E9, 1.666165545E9, 1.666165593E9, 1.666165641E9, 1.666165689E9, 1.666165737E9, 1.666165785E9, 1.666165833E9, 1.666165881E9, 1.666165929E9, 1.666165977E9, 1.666166025E9, 1.666166073E9, 1.666166121E9, 1.666166169E9, 1.66616652E9, 1.6661667E9, 1.66617052E9, 1.666170568E9, 1.666170616E9, 1.666170664E9, 1.666170712E9, 1.66617076E9, 1.666170808E9, 1.666170856E9, 1.666170904E9, 1.666170952E9, 1.666171E9, 1.666171048E9, 1.666171096E9, 1.666171144E9, 1.666171192E9, 1.66617124E9, 1.666171288E9, 1.666171336E9, 1.666171384E9, 1.666171432E9, 1.66617148E9, 1.666171528E9, 1.666171576E9, 1.666171624E9, 1.666171672E9, 1.66617172E9, 1.666171768E9, 1.666171816E9, 1.666171864E9, 1.666171912E9, 1.66617196E9, 1.666172008E9, 1.666172056E9, 1.666172104E9, 1.666172152E9, 1.6661722E9, 1.666172248E9, 1.666172296E9, 1.666172344E9, 1.666172392E9, 1.66617244E9, 1.6661727E9, 1.66617288E9, 1.666177362E9, 1.66617741E9, 1.666177458E9, 1.666177506E9, 1.666177554E9, 1.666177602E9, 1.66617765E9, 1.666177698E9, 1.666177746E9, 1.666177794E9, 1.666177842E9, 1.66617789E9, 1.666177938E9, 1.666177986E9, 1.666178034E9, 1.666178082E9, 1.66617813E9, 1.666178178E9, 1.666178226E9, 1.666178274E9, 1.666178322E9, 1.66617837E9, 1.666178418E9, 1.666178466E9, 1.666178514E9, 1.666178562E9, 1.66617861E9, 1.666178658E9, 1.666178706E9, 1.666178754E9, 1.666178802E9, 1.66617885E9, 1.666178898E9, 1.666178946E9, 1.666178994E9, 1.666179042E9, 1.66617909E9, 1.666179138E9, 1.666179186E9, 1.666179234E9, 1.666179282E9, 1.66617933E9, 1.666179378E9, 1.666179426E9, 1.666179474E9, 1.666179522E9, 1.66617957E9, 1.666179618E9, 1.666179666E9, 1.666179714E9, 1.666179762E9, 1.66617981E9, 1.66618008E9, 1.66618032E9, 1.666186219E9, 1.666186267E9, 1.666186315E9, 1.666186363E9, 1.666186411E9, 1.666186459E9, 1.666186507E9, 1.666186555E9, 1.666186603E9, 1.666186651E9, 1.666186699E9, 1.666186747E9, 1.666186795E9, 1.666186843E9, 1.666186891E9, 1.666186939E9, 1.666186987E9, 1.666187035E9, 1.666187083E9, 1.666187131E9, 1.666187179E9, 1.666187227E9, 1.666187275E9, 1.666187323E9, 1.666187371E9, 1.666187419E9, 1.666187467E9, 1.666187515E9, 1.666187563E9, 1.666187611E9, 1.666187659E9, 1.666187707E9, 1.666187755E9, 1.666187803E9, 1.666187851E9, 1.666187899E9, 1.666187947E9, 1.666187995E9, 1.666188043E9, 1.666188091E9, 1.666188139E9, 1.666188187E9, 1.666188235E9, 1.666188283E9, 1.666188331E9, 1.666188379E9, 1.666188427E9, 1.666188475E9, 1.666188523E9, 1.666188571E9, 1.666188619E9, 1.666188667E9, 1.666188715E9, 1.666188763E9, 1.666188811E9, 1.666188859E9, 1.666188907E9, 1.666188955E9, 1.666189003E9, 1.666189051E9, 1.666189099E9, 1.666189147E9, 1.666189195E9, 1.666189243E9, 1.666189291E9, 1.666189339E9, 1.666189387E9, 1.666189435E9, 1.666189483E9, 1.666189531E9, 1.666189579E9, 1.66618992E9, 1.66619016E9, 1.666195895E9, 1.666195943E9, 1.666195991E9, 1.666196039E9, 1.666196087E9, 1.666196135E9, 1.666196183E9, 1.666196231E9, 1.666196279E9, 1.666196327E9, 1.666196375E9, 1.666196423E9, 1.666196471E9, 1.666196519E9, 1.666196567E9, 1.666196615E9, 1.666196663E9, 1.666196711E9, 1.666196759E9, 1.666196807E9, 1.666196855E9, 1.666196903E9, 1.666196951E9, 1.666196999E9, 1.666197047E9, 1.666197095E9, 1.666197143E9, 1.666197191E9, 1.666197239E9, 1.666197287E9, 1.666197335E9, 1.666197383E9, 1.666197431E9, 1.666197479E9, 1.666197527E9, 1.666197575E9, 1.666197623E9, 1.666197671E9, 1.666197719E9, 1.666197767E9, 1.666197815E9, 1.666197863E9, 1.666197911E9, 1.666197959E9, 1.666198007E9, 1.666198055E9, 1.666198103E9, 1.666198151E9, 1.666198199E9, 1.666198247E9, 1.666198295E9, 1.666198343E9, 1.666198391E9, 1.666198439E9, 1.666198487E9, 1.666198535E9, 1.666198583E9, 1.666198631E9, 1.666198679E9, 1.666198727E9, 1.666198775E9, 1.666198823E9, 1.666198871E9, 1.666198919E9, 1.666198967E9, 1.666199015E9, 1.666199063E9, 1.666199111E9, 1.666199159E9, 1.66619958E9, 1.66619976E9, 1.666205612E9, 1.66620566E9, 1.666205708E9, 1.666205756E9, 1.666205804E9, 1.666205852E9, 1.6662059E9, 1.666205948E9, 1.666205996E9, 1.666206044E9, 1.666206092E9, 1.66620614E9, 1.666206188E9, 1.666206236E9, 1.666206284E9, 1.666206332E9, 1.66620638E9, 1.666206428E9, 1.666206476E9, 1.666206524E9, 1.666206572E9, 1.66620662E9, 1.666206668E9, 1.666206716E9, 1.666206764E9, 1.666206812E9, 1.66620686E9, 1.666206908E9, 1.666206956E9, 1.666207004E9, 1.666207052E9, 1.6662071E9, 1.666207148E9, 1.666207196E9, 1.666207244E9, 1.666207292E9, 1.66620734E9, 1.666207388E9, 1.666207436E9, 1.666207484E9, 1.666207532E9, 1.66620758E9, 1.666207628E9, 1.666207676E9, 1.666207724E9, 1.666207772E9, 1.66620782E9, 1.666207868E9, 1.666207916E9, 1.666207964E9, 1.666208012E9, 1.66620806E9, 1.666208108E9, 1.666208156E9, 1.666208204E9, 1.666208252E9, 1.6662083E9, 1.666208348E9, 1.666208396E9, 1.666208444E9, 1.666208492E9, 1.66620854E9, 1.666208588E9, 1.666208636E9, 1.666208684E9, 1.666208732E9, 1.66620878E9, 1.666208828E9, 1.666208876E9, 1.666208924E9, 1.666208972E9, 1.66620902E9, 1.6662093E9, 1.66620948E9, 1.666215372E9, 1.66621542E9, 1.666215468E9, 1.666215516E9, 1.666215564E9, 1.666215612E9, 1.66621566E9, 1.666215708E9, 1.666215756E9, 1.666215804E9, 1.666215852E9, 1.6662159E9, 1.666215948E9, 1.666215996E9, 1.666216044E9, 1.666216092E9, 1.66621614E9, 1.666216188E9, 1.666216236E9, 1.666216284E9, 1.666216332E9, 1.66621638E9, 1.666216428E9, 1.666216476E9, 1.666216524E9, 1.666216572E9, 1.66621662E9, 1.666216668E9, 1.666216716E9, 1.666216764E9, 1.666216812E9, 1.66621686E9, 1.666216908E9, 1.666216956E9, 1.666217004E9, 1.666217052E9, 1.6662171E9, 1.666217148E9, 1.666217196E9, 1.666217244E9, 1.666217292E9, 1.66621734E9, 1.666217388E9, 1.666217436E9, 1.666217484E9, 1.666217532E9, 1.66621758E9, 1.666217628E9, 1.666217676E9, 1.666217724E9, 1.666217772E9, 1.66621782E9, 1.666217868E9, 1.666217916E9, 1.666217964E9, 1.666218012E9, 1.66621806E9, 1.666218108E9, 1.666218156E9, 1.666218204E9, 1.666218252E9, 1.6662183E9, 1.666218348E9, 1.666218396E9, 1.666218444E9, 1.666218492E9, 1.66621854E9, 1.666218588E9, 1.666218636E9, 1.666218684E9, 1.666218732E9, 1.66621878E9, 1.6662192E9, 1.66621938E9, 1.666225242E9, 1.66622529E9, 1.666225338E9, 1.666225386E9, 1.666225434E9, 1.666225482E9, 1.66622553E9, 1.666225578E9, 1.666225626E9, 1.666225674E9, 1.666225722E9, 1.66622577E9, 1.666225818E9, 1.666225866E9, 1.666225914E9, 1.666225962E9, 1.66622601E9, 1.666226058E9, 1.666226106E9, 1.666226154E9, 1.666226202E9, 1.66622625E9, 1.666226298E9, 1.666226346E9, 1.666226394E9, 1.666226442E9, 1.66622649E9, 1.666226538E9, 1.666226586E9, 1.666226634E9, 1.666226682E9, 1.66622673E9, 1.666226778E9, 1.666226826E9, 1.666226874E9, 1.666226922E9, 1.66622697E9, 1.666227018E9, 1.666227066E9, 1.666227114E9, 1.666227162E9, 1.66622721E9, 1.666227258E9, 1.666227306E9, 1.666227354E9, 1.666227402E9, 1.66622745E9, 1.666227498E9, 1.666227546E9, 1.666227594E9, 1.666227642E9, 1.66622769E9, 1.666227738E9, 1.666227786E9, 1.666227834E9, 1.666227882E9, 1.66622793E9, 1.666227978E9, 1.666228026E9, 1.666228074E9, 1.666228122E9, 1.66622817E9, 1.666228218E9, 1.666228266E9, 1.666228314E9, 1.666228362E9, 1.66622841E9, 1.666228458E9, 1.666228506E9, 1.666228554E9, 1.666228602E9, 1.66622865E9, 1.66622898E9, 1.66622916E9, 1.666234999E9, 1.666235047E9, 1.666235095E9, 1.666235143E9, 1.666235191E9, 1.666235239E9, 1.666235287E9, 1.666235335E9, 1.666235383E9, 1.666235431E9, 1.666235479E9, 1.666235527E9, 1.666235575E9, 1.666235623E9, 1.666235671E9, 1.666235719E9, 1.666235767E9, 1.666235815E9, 1.666235863E9, 1.666235911E9, 1.666235959E9, 1.666236007E9, 1.666236055E9, 1.666236103E9, 1.666236151E9, 1.666236199E9, 1.666236247E9, 1.666236295E9, 1.666236343E9, 1.666236391E9, 1.666236439E9, 1.666236487E9, 1.666236535E9, 1.666236583E9, 1.666236631E9, 1.666236679E9, 1.666236727E9, 1.666236775E9, 1.666236823E9, 1.666236871E9, 1.666236919E9, 1.666236967E9, 1.666237015E9, 1.666237063E9, 1.666237111E9, 1.666237159E9, 1.666237207E9, 1.666237255E9, 1.666237303E9, 1.666237351E9, 1.666237399E9, 1.666237447E9, 1.666237495E9, 1.666237543E9, 1.666237591E9, 1.666237639E9, 1.666237687E9, 1.666237735E9, 1.666237783E9, 1.666237831E9, 1.666237879E9, 1.666237927E9, 1.666237975E9, 1.666238023E9, 1.666238071E9, 1.666238119E9, 1.666238167E9, 1.666238215E9, 1.666238263E9, 1.666238311E9, 1.666238359E9, 1.6662387E9, 1.66623888E9, 1.666244728E9, 1.666244776E9, 1.666244824E9, 1.666244872E9, 1.66624492E9, 1.666244968E9, 1.666245016E9, 1.666245064E9, 1.666245112E9, 1.66624516E9, 1.666245208E9, 1.666245256E9, 1.666245304E9, 1.666245352E9, 1.6662454E9, 1.666245448E9, 1.666245496E9, 1.666245544E9, 1.666245592E9, 1.66624564E9, 1.666245688E9, 1.666245736E9, 1.666245784E9, 1.666245832E9, 1.66624588E9, 1.666245928E9, 1.666245976E9, 1.666246024E9, 1.666246072E9, 1.66624612E9, 1.666246168E9, 1.666246216E9, 1.666246264E9, 1.666246312E9, 1.66624636E9, 1.666246408E9, 1.666246456E9, 1.666246504E9, 1.666246552E9, 1.6662466E9, 1.666246648E9, 1.666246696E9, 1.666246744E9, 1.666246792E9, 1.66624684E9, 1.666246888E9, 1.666246936E9, 1.666246984E9, 1.666247032E9, 1.66624708E9, 1.666247128E9, 1.666247176E9, 1.666247224E9, 1.666247272E9, 1.66624732E9, 1.666247368E9, 1.666247416E9, 1.666247464E9, 1.666247512E9, 1.66624756E9, 1.666247608E9, 1.666247656E9, 1.666247704E9, 1.666247752E9, 1.6662478E9, 1.666247848E9, 1.666247896E9, 1.666247944E9, 1.666247992E9, 1.66624804E9, 1.66624842E9, 1.6662486E9, 1.666254506E9, 1.666254554E9, 1.666254602E9, 1.66625465E9, 1.666254698E9, 1.666254746E9, 1.666254794E9, 1.666254842E9, 1.66625489E9, 1.666254938E9, 1.666254986E9, 1.666255034E9, 1.666255082E9, 1.66625513E9, 1.666255178E9, 1.666255226E9, 1.666255274E9, 1.666255322E9, 1.66625537E9, 1.666255418E9, 1.666255466E9, 1.666255514E9, 1.666255562E9, 1.66625561E9, 1.666255658E9, 1.666255706E9, 1.666255754E9, 1.666255802E9, 1.66625585E9, 1.666255898E9, 1.666255946E9, 1.666255994E9, 1.666256042E9, 1.66625609E9, 1.666256138E9, 1.666256186E9, 1.666256234E9, 1.666256282E9, 1.66625633E9, 1.666256378E9, 1.666256426E9, 1.666256474E9, 1.666256522E9, 1.66625657E9, 1.666256618E9, 1.666256666E9, 1.666256714E9, 1.666256762E9, 1.66625681E9, 1.666256858E9, 1.666256906E9, 1.666256954E9, 1.666257002E9, 1.66625705E9, 1.666257098E9, 1.666257146E9, 1.666257194E9, 1.666257242E9, 1.66625729E9, 1.666257338E9, 1.666257386E9, 1.666257434E9, 1.666257482E9, 1.66625753E9, 1.666257578E9, 1.666257626E9, 1.666257674E9, 1.666257722E9, 1.66625777E9, 1.666257818E9, 1.666257866E9, 1.666257914E9, 1.666257962E9, 1.66625801E9, 1.66625838E9, 1.66625856E9, 1.666264393E9, 1.666264441E9, 1.666264489E9, 1.666264537E9, 1.666264585E9, 1.666264633E9, 1.666264681E9, 1.666264729E9, 1.666264777E9, 1.666264825E9, 1.666264873E9, 1.666264921E9, 1.666264969E9, 1.666265017E9, 1.666265065E9, 1.666265113E9, 1.666265161E9, 1.666265209E9, 1.666265257E9, 1.666265305E9, 1.666265353E9, 1.666265401E9, 1.666265449E9, 1.666265497E9, 1.666265545E9, 1.666265593E9, 1.666265641E9, 1.666265689E9, 1.666265737E9, 1.666265785E9, 1.666265833E9, 1.666265881E9, 1.666265929E9, 1.666265977E9, 1.666266025E9, 1.666266073E9, 1.666266121E9, 1.666266169E9, 1.666266217E9, 1.666266265E9, 1.666266313E9, 1.666266361E9, 1.666266409E9, 1.666266457E9, 1.666266505E9, 1.666266553E9, 1.666266601E9, 1.666266649E9, 1.666266697E9, 1.666266745E9, 1.666266793E9, 1.666266841E9, 1.666266889E9, 1.666266937E9, 1.666266985E9, 1.666267033E9, 1.666267081E9, 1.666267129E9, 1.666267177E9, 1.666267225E9, 1.666267273E9, 1.666267321E9, 1.666267369E9, 1.666267417E9, 1.666267465E9, 1.666267513E9, 1.666267561E9, 1.666267609E9, 1.666267657E9, 1.666267705E9, 1.666267753E9, 1.666267801E9, 1.666267849E9, 1.666267897E9, 1.666267945E9, 1.666267993E9, 1.666268041E9, 1.666268089E9, 1.66626846E9, 1.66626864E9, 1.666274399E9, 1.666274447E9, 1.666274495E9, 1.666274543E9, 1.666274591E9, 1.666274639E9, 1.666274687E9, 1.666274735E9, 1.666274783E9, 1.666274831E9, 1.666274879E9, 1.666274927E9, 1.666274975E9, 1.666275023E9, 1.666275071E9, 1.666275119E9, 1.666275167E9, 1.666275215E9, 1.666275263E9, 1.666275311E9, 1.666275359E9, 1.666275407E9, 1.666275455E9, 1.666275503E9, 1.666275551E9, 1.666275599E9, 1.666275647E9, 1.666275695E9, 1.666275743E9, 1.666275791E9, 1.666275839E9, 1.666275887E9, 1.666275935E9, 1.666275983E9, 1.666276031E9, 1.666276079E9, 1.666276127E9, 1.666276175E9, 1.666276223E9, 1.666276271E9, 1.666276319E9, 1.666276367E9, 1.666276415E9, 1.666276463E9, 1.666276511E9, 1.666276559E9, 1.666276607E9, 1.666276655E9, 1.666276703E9, 1.666276751E9, 1.666276799E9, 1.666276847E9, 1.666276895E9, 1.666276943E9, 1.666276991E9, 1.666277039E9, 1.666277087E9, 1.666277135E9, 1.666277183E9, 1.666277231E9, 1.666277279E9, 1.666277327E9, 1.666277375E9, 1.666277423E9, 1.666277471E9, 1.666277519E9, 1.666277567E9, 1.666277615E9, 1.666277663E9, 1.666277711E9, 1.666277759E9, 1.666277807E9, 1.666277855E9, 1.666277903E9, 1.666277951E9, 1.666277999E9, 1.66627836E9, 1.66627854E9, 1.666284272E9, 1.66628432E9, 1.666284368E9, 1.666284416E9, 1.666284464E9, 1.666284512E9, 1.66628456E9, 1.666284608E9, 1.666284656E9, 1.666284704E9, 1.666284752E9, 1.6662848E9, 1.666284848E9, 1.666284896E9, 1.666284944E9, 1.666284992E9, 1.66628504E9, 1.666285088E9, 1.666285136E9, 1.666285184E9, 1.666285232E9, 1.66628528E9, 1.666285328E9, 1.666285376E9, 1.666285424E9, 1.666285472E9, 1.66628552E9, 1.666285568E9, 1.666285616E9, 1.666285664E9, 1.666285712E9, 1.66628576E9, 1.666285808E9, 1.666285856E9, 1.666285904E9, 1.666285952E9, 1.666286E9, 1.666286048E9, 1.666286096E9, 1.666286144E9, 1.666286192E9, 1.66628624E9, 1.666286288E9, 1.666286336E9, 1.666286384E9, 1.666286432E9, 1.66628648E9, 1.666286528E9, 1.666286576E9, 1.666286624E9, 1.666286672E9, 1.66628672E9, 1.666286768E9, 1.666286816E9, 1.666286864E9, 1.666286912E9, 1.66628696E9, 1.666287008E9, 1.666287056E9, 1.666287104E9, 1.666287152E9, 1.6662872E9, 1.666287248E9, 1.666287296E9, 1.666287344E9, 1.666287392E9, 1.66628744E9, 1.666287488E9, 1.666287536E9, 1.666287584E9, 1.666287632E9, 1.66628768E9, 1.66628808E9, 1.66628826E9, 1.666293912E9, 1.66629396E9, 1.666294008E9, 1.666294056E9, 1.666294104E9, 1.666294152E9, 1.6662942E9, 1.666294248E9, 1.666294296E9, 1.666294344E9, 1.666294392E9, 1.66629444E9, 1.666294488E9, 1.666294536E9, 1.666294584E9, 1.666294632E9, 1.66629468E9, 1.666294728E9, 1.666294776E9, 1.666294824E9, 1.666294872E9, 1.66629492E9, 1.666294968E9, 1.666295016E9, 1.666295064E9, 1.666295112E9, 1.66629516E9, 1.666295208E9, 1.666295256E9, 1.666295304E9, 1.666295352E9, 1.6662954E9, 1.666295448E9, 1.666295496E9, 1.666295544E9, 1.666295592E9, 1.66629564E9, 1.666295688E9, 1.666295736E9, 1.666295784E9, 1.666295832E9, 1.66629588E9, 1.666295928E9, 1.666295976E9, 1.666296024E9, 1.666296072E9, 1.66629612E9, 1.666296168E9, 1.666296216E9, 1.666296264E9, 1.666296312E9, 1.66629636E9, 1.666296408E9, 1.666296456E9, 1.666296504E9, 1.666296552E9, 1.6662966E9, 1.666296648E9, 1.666296696E9, 1.666296744E9, 1.666296792E9, 1.66629684E9, 1.666296888E9, 1.666296936E9, 1.666296984E9, 1.666297032E9, 1.66629708E9, 1.666297128E9, 1.666297176E9, 1.666297224E9, 1.666297272E9, 1.66629732E9, 1.66629774E9, 1.66629798E9, 1.666303772E9, 1.66630382E9, 1.666303868E9, 1.666303916E9, 1.666303964E9, 1.666304012E9, 1.66630406E9, 1.666304108E9, 1.666304156E9, 1.666304204E9, 1.666304252E9, 1.6663043E9, 1.666304348E9, 1.666304396E9, 1.666304444E9, 1.666304492E9, 1.66630454E9, 1.666304588E9, 1.666304636E9, 1.666304684E9, 1.666304732E9, 1.66630478E9, 1.666304828E9, 1.666304876E9, 1.666304924E9, 1.666304972E9, 1.66630502E9, 1.666305068E9, 1.666305116E9, 1.666305164E9, 1.666305212E9, 1.66630526E9, 1.666305308E9, 1.666305356E9, 1.666305404E9, 1.666305452E9, 1.6663055E9, 1.666305548E9, 1.666305596E9, 1.666305644E9, 1.666305692E9, 1.66630574E9, 1.666305788E9, 1.666305836E9, 1.666305884E9, 1.666305932E9, 1.66630598E9, 1.666306028E9, 1.666306076E9, 1.666306124E9, 1.666306172E9, 1.66630622E9, 1.666306268E9, 1.666306316E9, 1.666306364E9, 1.666306412E9, 1.66630646E9, 1.666306508E9, 1.666306556E9, 1.666306604E9, 1.666306652E9, 1.6663067E9, 1.666306748E9, 1.666306796E9, 1.666306844E9, 1.666306892E9, 1.66630694E9, 1.666306988E9, 1.666307036E9, 1.666307084E9, 1.666307132E9, 1.66630718E9, 1.66630752E9, 1.6663077E9, 1.666313416E9, 1.666313464E9, 1.666313512E9, 1.66631356E9, 1.666313608E9, 1.666313656E9, 1.666313704E9, 1.666313752E9, 1.6663138E9, 1.666313848E9, 1.666313896E9, 1.666313944E9, 1.666313992E9, 1.66631404E9, 1.666314088E9, 1.666314136E9, 1.666314184E9, 1.666314232E9, 1.66631428E9, 1.666314328E9, 1.666314376E9, 1.666314424E9, 1.666314472E9, 1.66631452E9, 1.666314568E9, 1.666314616E9, 1.666314664E9, 1.666314712E9, 1.66631476E9, 1.666314808E9, 1.666314856E9, 1.666314904E9, 1.666314952E9, 1.666315E9, 1.666315048E9, 1.666315096E9, 1.666315144E9, 1.666315192E9, 1.66631524E9, 1.666315288E9, 1.666315336E9, 1.666315384E9, 1.666315432E9, 1.66631548E9, 1.666315528E9, 1.666315576E9, 1.666315624E9, 1.666315672E9, 1.66631572E9, 1.666315768E9, 1.666315816E9, 1.666315864E9, 1.666315912E9, 1.66631596E9, 1.666316008E9, 1.666316056E9, 1.666316104E9, 1.666316152E9, 1.6663162E9, 1.666316248E9, 1.666316296E9, 1.666316344E9, 1.666316392E9, 1.66631644E9, 1.666316488E9, 1.666316536E9, 1.666316584E9, 1.666316632E9, 1.66631668E9, 1.666316728E9, 1.666316776E9, 1.666316824E9, 1.666316872E9, 1.66631692E9, 1.6663173E9, 1.66631742E9, 1.666323395E9, 1.666323443E9, 1.666323491E9, 1.666323539E9, 1.666323587E9, 1.666323635E9, 1.666323683E9, 1.666323731E9, 1.666323779E9, 1.666323827E9, 1.666323875E9, 1.666323923E9, 1.666323971E9, 1.666324019E9, 1.666324067E9, 1.666324115E9, 1.666324163E9, 1.666324211E9, 1.666324259E9, 1.666324307E9, 1.666324355E9, 1.666324403E9, 1.666324451E9, 1.666324499E9, 1.666324547E9, 1.666324595E9, 1.666324643E9, 1.666324691E9, 1.666324739E9, 1.666324787E9, 1.666324835E9, 1.666324883E9, 1.666324931E9, 1.666324979E9, 1.666325027E9, 1.666325075E9, 1.666325123E9, 1.666325171E9, 1.666325219E9, 1.666325267E9, 1.666325315E9, 1.666325363E9, 1.666325411E9, 1.666325459E9, 1.666325507E9, 1.666325555E9, 1.666325603E9, 1.666325651E9, 1.666325699E9, 1.666325747E9, 1.666325795E9, 1.666325843E9, 1.666325891E9, 1.666325939E9, 1.666325987E9, 1.666326035E9, 1.666326083E9, 1.666326131E9, 1.666326179E9, 1.666326227E9, 1.666326275E9, 1.666326323E9, 1.666326371E9, 1.666326419E9, 1.666326467E9, 1.666326515E9, 1.666326563E9, 1.666326611E9, 1.666326659E9, 1.666326707E9, 1.666326755E9, 1.666326803E9, 1.666326851E9, 1.666326899E9, 1.66632732E9, 1.666327321E9, 1.66633339E9, 1.666333438E9, 1.666333486E9, 1.666333534E9, 1.666333582E9, 1.66633363E9, 1.666333678E9, 1.666333726E9, 1.666333774E9, 1.666333822E9, 1.66633387E9, 1.666333918E9, 1.666333966E9, 1.666334014E9, 1.666334062E9, 1.66633411E9, 1.666334158E9, 1.666334206E9, 1.666334254E9, 1.666334302E9, 1.66633435E9, 1.666334398E9, 1.666334446E9, 1.666334494E9, 1.666334542E9, 1.66633459E9, 1.666334638E9, 1.666334686E9, 1.666334734E9, 1.666334782E9, 1.66633483E9, 1.666334878E9, 1.666334926E9, 1.666334974E9, 1.666335022E9, 1.66633507E9, 1.666335118E9, 1.666335166E9, 1.666335214E9, 1.666335262E9, 1.66633531E9, 1.666335358E9, 1.666335406E9, 1.666335454E9, 1.666335502E9, 1.66633555E9, 1.666335598E9, 1.666335646E9, 1.666335694E9, 1.666335742E9, 1.66633579E9, 1.666335838E9, 1.666335886E9, 1.666335934E9, 1.666335982E9, 1.66633603E9, 1.666336078E9, 1.666336126E9, 1.666336174E9, 1.666336222E9, 1.66633627E9, 1.666336318E9, 1.666336366E9, 1.666336414E9, 1.666336462E9, 1.66633651E9, 1.666336558E9, 1.666336606E9, 1.666336654E9, 1.666336702E9, 1.66633675E9, 1.66633716E9, 1.666337161E9, 1.666342819E9, 1.666342867E9, 1.666342915E9, 1.666342963E9, 1.666343011E9, 1.666343059E9, 1.666343107E9, 1.666343155E9, 1.666343203E9, 1.666343251E9, 1.666343299E9, 1.666343347E9, 1.666343395E9, 1.666343443E9, 1.666343491E9, 1.666343539E9, 1.666343587E9, 1.666343635E9, 1.666343683E9, 1.666343731E9, 1.666343779E9, 1.666343827E9, 1.666343875E9, 1.666343923E9, 1.666343971E9, 1.666344019E9, 1.666344067E9, 1.666344115E9, 1.666344163E9, 1.666344211E9, 1.666344259E9, 1.666344307E9, 1.666344355E9, 1.666344403E9, 1.666344451E9, 1.666344499E9, 1.666344547E9, 1.666344595E9, 1.666344643E9, 1.666344691E9, 1.666344739E9, 1.666344787E9, 1.666344835E9, 1.666344883E9, 1.666344931E9, 1.666344979E9, 1.666345027E9, 1.666345075E9, 1.666345123E9, 1.666345171E9, 1.666345219E9, 1.666345267E9, 1.666345315E9, 1.666345363E9, 1.666345411E9, 1.666345459E9, 1.666345507E9, 1.666345555E9, 1.666345603E9, 1.666345651E9, 1.666345699E9, 1.666345747E9, 1.666345795E9, 1.666345843E9, 1.666345891E9, 1.666345939E9, 1.666345987E9, 1.666346035E9, 1.666346083E9, 1.666346131E9, 1.666346179E9, 1.66634658E9, 1.66634676E9, 1.66635243E9, 1.666352478E9, 1.666352526E9, 1.666352574E9, 1.666352622E9, 1.66635267E9, 1.666352718E9, 1.666352766E9, 1.666352814E9, 1.666352862E9, 1.66635291E9, 1.666352958E9, 1.666353006E9, 1.666353054E9, 1.666353102E9, 1.66635315E9, 1.666353198E9, 1.666353246E9, 1.666353294E9, 1.666353342E9, 1.66635339E9, 1.666353438E9, 1.666353486E9, 1.666353534E9, 1.666353582E9, 1.66635363E9, 1.666353678E9, 1.666353726E9, 1.666353774E9, 1.666353822E9, 1.66635387E9, 1.666353918E9, 1.666353966E9, 1.666354014E9, 1.666354062E9, 1.66635411E9, 1.666354158E9, 1.666354206E9, 1.666354254E9, 1.666354302E9, 1.66635435E9, 1.666354398E9, 1.666354446E9, 1.666354494E9, 1.666354542E9, 1.66635459E9, 1.666354638E9, 1.666354686E9, 1.666354734E9, 1.666354782E9, 1.66635483E9, 1.666354878E9, 1.666354926E9, 1.666354974E9, 1.666355022E9, 1.66635507E9, 1.666355118E9, 1.666355166E9, 1.666355214E9, 1.666355262E9, 1.66635531E9, 1.666355358E9, 1.666355406E9, 1.666355454E9, 1.666355502E9, 1.66635555E9, 1.666355598E9, 1.666355646E9, 1.666355694E9, 1.666355742E9, 1.66635579E9, 1.66635606E9, 1.6663563E9, 1.666361971E9, 1.666362019E9, 1.666362067E9, 1.666362115E9, 1.666362163E9, 1.666362211E9, 1.666362259E9, 1.666362307E9, 1.666362355E9, 1.666362403E9, 1.666362451E9, 1.666362499E9, 1.666362547E9, 1.666362595E9, 1.666362643E9, 1.666362691E9, 1.666362739E9, 1.666362787E9, 1.666362835E9, 1.666362883E9, 1.666362931E9, 1.666362979E9, 1.666363027E9, 1.666363075E9, 1.666363123E9, 1.666363171E9, 1.666363219E9, 1.666363267E9, 1.666363315E9, 1.666363363E9, 1.666363411E9, 1.666363459E9, 1.666363507E9, 1.666363555E9, 1.666363603E9, 1.666363651E9, 1.666363699E9, 1.666363747E9, 1.666363795E9, 1.666363843E9, 1.666363891E9, 1.666363939E9, 1.666363987E9, 1.666364035E9, 1.666364083E9, 1.666364131E9, 1.666364179E9, 1.666364227E9, 1.666364275E9, 1.666364323E9, 1.666364371E9, 1.666364419E9, 1.666364467E9, 1.666364515E9, 1.666364563E9, 1.666364611E9, 1.666364659E9, 1.666364707E9, 1.666364755E9, 1.666364803E9, 1.666364851E9, 1.666364899E9, 1.666364947E9, 1.666364995E9, 1.666365043E9, 1.666365091E9, 1.666365139E9, 1.666365187E9, 1.666365235E9, 1.666365283E9, 1.666365331E9, 1.666365379E9, 1.66636566E9, 1.6663659E9, 1.666371682E9, 1.66637173E9, 1.666371778E9, 1.666371826E9, 1.666371874E9, 1.666371922E9, 1.66637197E9, 1.666372018E9, 1.666372066E9, 1.666372114E9, 1.666372162E9, 1.66637221E9, 1.666372258E9, 1.666372306E9, 1.666372354E9, 1.666372402E9, 1.66637245E9, 1.666372498E9, 1.666372546E9, 1.666372594E9, 1.666372642E9, 1.66637269E9, 1.666372738E9, 1.666372786E9, 1.666372834E9, 1.666372882E9, 1.66637293E9, 1.666372978E9, 1.666373026E9, 1.666373074E9, 1.666373122E9, 1.66637317E9, 1.666373218E9, 1.666373266E9, 1.666373314E9, 1.666373362E9, 1.66637341E9, 1.666373458E9, 1.666373506E9, 1.666373554E9, 1.666373602E9, 1.66637365E9, 1.666373698E9, 1.666373746E9, 1.666373794E9, 1.666373842E9, 1.66637389E9, 1.666373938E9, 1.666373986E9, 1.666374034E9, 1.666374082E9, 1.66637413E9, 1.666374178E9, 1.666374226E9, 1.666374274E9, 1.666374322E9, 1.66637437E9, 1.666374418E9, 1.666374466E9, 1.666374514E9, 1.666374562E9, 1.66637461E9, 1.666374658E9, 1.666374706E9, 1.666374754E9, 1.666374802E9, 1.66637485E9, 1.666374898E9, 1.666374946E9, 1.666374994E9, 1.666375042E9, 1.66637509E9, 1.6663755E9, 1.66637568E9, 1.666381678E9, 1.666381726E9, 1.666381774E9, 1.666381822E9, 1.66638187E9, 1.666381918E9, 1.666381966E9, 1.666382014E9, 1.666382062E9, 1.66638211E9, 1.666382158E9, 1.666382206E9, 1.666382254E9, 1.666382302E9, 1.66638235E9, 1.666382398E9, 1.666382446E9, 1.666382494E9, 1.666382542E9, 1.66638259E9, 1.666382638E9, 1.666382686E9, 1.666382734E9, 1.666382782E9, 1.66638283E9, 1.666382878E9, 1.666382926E9, 1.666382974E9, 1.666383022E9, 1.66638307E9, 1.666383118E9, 1.666383166E9, 1.666383214E9, 1.666383262E9, 1.66638331E9, 1.666383358E9, 1.666383406E9, 1.666383454E9, 1.666383502E9, 1.66638355E9, 1.666383598E9, 1.666383646E9, 1.666383694E9, 1.666383742E9, 1.66638379E9, 1.666383838E9, 1.666383886E9, 1.666383934E9, 1.666383982E9, 1.66638403E9, 1.666384078E9, 1.666384126E9, 1.666384174E9, 1.666384222E9, 1.66638427E9, 1.666384318E9, 1.666384366E9, 1.666384414E9, 1.666384462E9, 1.66638451E9, 1.666384558E9, 1.666384606E9, 1.666384654E9, 1.666384702E9, 1.66638475E9, 1.666384798E9, 1.666384846E9, 1.666384894E9, 1.666384942E9, 1.66638499E9, 1.66638528E9, 1.66638546E9, 1.666391368E9, 1.666391416E9, 1.666391464E9, 1.666391512E9, 1.66639156E9, 1.666391608E9, 1.666391656E9, 1.666391704E9, 1.666391752E9, 1.6663918E9, 1.666391848E9, 1.666391896E9, 1.666391944E9, 1.666391992E9, 1.66639204E9, 1.666392088E9, 1.666392136E9, 1.666392184E9, 1.666392232E9, 1.66639228E9, 1.666392328E9, 1.666392376E9, 1.666392424E9, 1.666392472E9, 1.66639252E9, 1.666392568E9, 1.666392616E9, 1.666392664E9, 1.666392712E9, 1.66639276E9, 1.666392808E9, 1.666392856E9, 1.666392904E9, 1.666392952E9, 1.666393E9, 1.666393048E9, 1.666393096E9, 1.666393144E9, 1.666393192E9, 1.66639324E9, 1.666393288E9, 1.666393336E9, 1.666393384E9, 1.666393432E9, 1.66639348E9, 1.666393528E9, 1.666393576E9, 1.666393624E9, 1.666393672E9, 1.66639372E9, 1.666393768E9, 1.666393816E9, 1.666393864E9, 1.666393912E9, 1.66639396E9, 1.666394008E9, 1.666394056E9, 1.666394104E9, 1.666394152E9, 1.6663942E9, 1.666394248E9, 1.666394296E9, 1.666394344E9, 1.666394392E9, 1.66639444E9, 1.666394488E9, 1.666394536E9, 1.666394584E9, 1.666394632E9, 1.66639468E9, 1.666394728E9, 1.666394776E9, 1.666394824E9, 1.666394872E9, 1.66639492E9, 1.66639524E9, 1.66639542E9, 1.666401046E9, 1.666401094E9, 1.666401142E9, 1.66640119E9, 1.666401238E9, 1.666401286E9, 1.666401334E9, 1.666401382E9, 1.66640143E9, 1.666401478E9, 1.666401526E9, 1.666401574E9, 1.666401622E9, 1.66640167E9, 1.666401718E9, 1.666401766E9, 1.666401814E9, 1.666401862E9, 1.66640191E9, 1.666401958E9, 1.666402006E9, 1.666402054E9, 1.666402102E9, 1.66640215E9, 1.666402198E9, 1.666402246E9, 1.666402294E9, 1.666402342E9, 1.66640239E9, 1.666402438E9, 1.666402486E9, 1.666402534E9, 1.666402582E9, 1.66640263E9, 1.666402678E9, 1.666402726E9, 1.666402774E9, 1.666402822E9, 1.66640287E9, 1.666402918E9, 1.666402966E9, 1.666403014E9, 1.666403062E9, 1.66640311E9, 1.666403158E9, 1.666403206E9, 1.666403254E9, 1.666403302E9, 1.66640335E9, 1.666403398E9, 1.666403446E9, 1.666403494E9, 1.666403542E9, 1.66640359E9, 1.666403638E9, 1.666403686E9, 1.666403734E9, 1.666403782E9, 1.66640383E9, 1.666403878E9, 1.666403926E9, 1.666403974E9, 1.666404022E9, 1.66640407E9, 1.666404118E9, 1.666404166E9, 1.666404214E9, 1.666404262E9, 1.66640431E9, 1.66640472E9, 1.6664049E9, 1.666410924E9, 1.666410972E9, 1.66641102E9, 1.666411068E9, 1.666411116E9, 1.666411164E9, 1.666411212E9, 1.66641126E9, 1.666411308E9, 1.666411356E9, 1.666411404E9, 1.666411452E9, 1.6664115E9, 1.666411548E9, 1.666411596E9, 1.666411644E9, 1.666411692E9, 1.66641174E9, 1.666411788E9, 1.666411836E9, 1.666411884E9, 1.666411932E9, 1.66641198E9, 1.666412028E9, 1.666412076E9, 1.666412124E9, 1.666412172E9, 1.66641222E9, 1.666412268E9, 1.666412316E9, 1.666412364E9, 1.666412412E9, 1.66641246E9, 1.666412508E9, 1.666412556E9, 1.666412604E9, 1.666412652E9, 1.6664127E9, 1.666412748E9, 1.666412796E9, 1.666412844E9, 1.666412892E9, 1.66641294E9, 1.666412988E9, 1.666413036E9, 1.666413084E9, 1.666413132E9, 1.66641318E9, 1.666413228E9, 1.666413276E9, 1.666413324E9, 1.666413372E9, 1.66641342E9, 1.666413468E9, 1.666413516E9, 1.666413564E9, 1.666413612E9, 1.66641366E9, 1.666413708E9, 1.666413756E9, 1.666413804E9, 1.666413852E9, 1.6664139E9, 1.666413948E9, 1.666413996E9, 1.666414044E9, 1.666414092E9, 1.66641414E9, 1.666414188E9, 1.666414236E9, 1.666414284E9, 1.666414332E9, 1.66641438E9, 1.6664148E9, 1.666414801E9, 1.666420596E9, 1.666420644E9, 1.666420692E9, 1.66642074E9, 1.666420788E9, 1.666420836E9, 1.666420884E9, 1.666420932E9, 1.66642098E9, 1.666421028E9, 1.666421076E9, 1.666421124E9, 1.666421172E9, 1.66642122E9, 1.666421268E9, 1.666421316E9, 1.666421364E9, 1.666421412E9, 1.66642146E9, 1.666421508E9, 1.666421556E9, 1.666421604E9, 1.666421652E9, 1.6664217E9, 1.666421748E9, 1.666421796E9, 1.666421844E9, 1.666421892E9, 1.66642194E9, 1.666421988E9, 1.666422036E9, 1.666422084E9, 1.666422132E9, 1.66642218E9, 1.666422228E9, 1.666422276E9, 1.666422324E9, 1.666422372E9, 1.66642242E9, 1.666422468E9, 1.666422516E9, 1.666422564E9, 1.666422612E9, 1.66642266E9, 1.666422708E9, 1.666422756E9, 1.666422804E9, 1.666422852E9, 1.6664229E9, 1.666422948E9, 1.666422996E9, 1.666423044E9, 1.666423092E9, 1.66642314E9, 1.666423188E9, 1.666423236E9, 1.666423284E9, 1.666423332E9, 1.66642338E9, 1.666423428E9, 1.666423476E9, 1.666423524E9, 1.666423572E9, 1.66642362E9, 1.666423668E9, 1.666423716E9, 1.666423764E9, 1.666423812E9, 1.66642386E9, 1.666423908E9, 1.666423956E9, 1.666424004E9, 1.666424052E9, 1.6664241E9, 1.6664244E9, 1.66642464E9, 1.666430392E9, 1.66643044E9, 1.666430488E9, 1.666430536E9, 1.666430584E9, 1.666430632E9, 1.66643068E9, 1.666430728E9, 1.666430776E9, 1.666430824E9, 1.666430872E9, 1.66643092E9, 1.666430968E9, 1.666431016E9, 1.666431064E9, 1.666431112E9, 1.66643116E9, 1.666431208E9, 1.666431256E9, 1.666431304E9, 1.666431352E9, 1.6664314E9, 1.666431448E9, 1.666431496E9, 1.666431544E9, 1.666431592E9, 1.66643164E9, 1.666431688E9, 1.666431736E9, 1.666431784E9, 1.666431832E9, 1.66643188E9, 1.666431928E9, 1.666431976E9, 1.666432024E9, 1.666432072E9, 1.66643212E9, 1.666432168E9, 1.666432216E9, 1.666432264E9, 1.666432312E9, 1.66643236E9, 1.666432408E9, 1.666432456E9, 1.666432504E9, 1.666432552E9, 1.6664326E9, 1.666432648E9, 1.666432696E9, 1.666432744E9, 1.666432792E9, 1.66643284E9, 1.666432888E9, 1.666432936E9, 1.666432984E9, 1.666433032E9, 1.66643308E9, 1.666433128E9, 1.666433176E9, 1.666433224E9, 1.666433272E9, 1.66643332E9, 1.666433368E9, 1.666433416E9, 1.666433464E9, 1.666433512E9, 1.66643356E9, 1.666433608E9, 1.666433656E9, 1.666433704E9, 1.666433752E9, 1.6664338E9, 1.66643418E9, 1.66643436E9, 1.666440105E9, 1.666440153E9, 1.666440201E9, 1.666440249E9, 1.666440297E9, 1.666440345E9, 1.666440393E9, 1.666440441E9, 1.666440489E9, 1.666440537E9, 1.666440585E9, 1.666440633E9, 1.666440681E9, 1.666440729E9, 1.666440777E9, 1.666440825E9, 1.666440873E9, 1.666440921E9, 1.666440969E9, 1.666441017E9, 1.666441065E9, 1.666441113E9, 1.666441161E9, 1.666441209E9, 1.666441257E9, 1.666441305E9, 1.666441353E9, 1.666441401E9, 1.666441449E9, 1.666441497E9, 1.666441545E9, 1.666441593E9, 1.666441641E9, 1.666441689E9, 1.666441737E9, 1.666441785E9, 1.666441833E9, 1.666441881E9, 1.666441929E9, 1.666441977E9, 1.666442025E9, 1.666442073E9, 1.666442121E9, 1.666442169E9, 1.666442217E9, 1.666442265E9, 1.666442313E9, 1.666442361E9, 1.666442409E9, 1.666442457E9, 1.666442505E9, 1.666442553E9, 1.666442601E9, 1.666442649E9, 1.666442697E9, 1.666442745E9, 1.666442793E9, 1.666442841E9, 1.666442889E9, 1.666442937E9, 1.666442985E9, 1.666443033E9, 1.666443081E9, 1.666443129E9, 1.666443177E9, 1.666443225E9, 1.666443273E9, 1.666443321E9, 1.666443369E9, 1.66644378E9, 1.66644396E9, 1.666449587E9, 1.666449635E9, 1.666449683E9, 1.666449731E9, 1.666449779E9, 1.666449827E9, 1.666449875E9, 1.666449923E9, 1.666449971E9, 1.666450019E9, 1.666450067E9, 1.666450115E9, 1.666450163E9, 1.666450211E9, 1.666450259E9, 1.666450307E9, 1.666450355E9, 1.666450403E9, 1.666450451E9, 1.666450499E9, 1.666450547E9, 1.666450595E9, 1.666450643E9, 1.666450691E9, 1.666450739E9, 1.666450787E9, 1.666450835E9, 1.666450883E9, 1.666450931E9, 1.666450979E9, 1.666451027E9, 1.666451075E9, 1.666451123E9, 1.666451171E9, 1.666451219E9, 1.666451267E9, 1.666451315E9, 1.666451363E9, 1.666451411E9, 1.666451459E9, 1.666451507E9, 1.666451555E9, 1.666451603E9, 1.666451651E9, 1.666451699E9, 1.666451747E9, 1.666451795E9, 1.666451843E9, 1.666451891E9, 1.666451939E9, 1.666451987E9, 1.666452035E9, 1.666452083E9, 1.666452131E9, 1.666452179E9, 1.666452227E9, 1.666452275E9, 1.666452323E9, 1.666452371E9, 1.666452419E9, 1.666452467E9, 1.666452515E9, 1.666452563E9, 1.666452611E9, 1.666452659E9, 1.666452707E9, 1.666452755E9, 1.666452803E9, 1.666452851E9, 1.666452899E9, 1.6664532E9, 1.66645338E9, 1.666459338E9, 1.666459386E9, 1.666459434E9, 1.666459482E9, 1.66645953E9, 1.666459578E9, 1.666459626E9, 1.666459674E9, 1.666459722E9, 1.66645977E9, 1.666459818E9, 1.666459866E9, 1.666459914E9, 1.666459962E9, 1.66646001E9, 1.666460058E9, 1.666460106E9, 1.666460154E9, 1.666460202E9, 1.66646025E9, 1.666460298E9, 1.666460346E9, 1.666460394E9, 1.666460442E9, 1.66646049E9, 1.666460538E9, 1.666460586E9, 1.666460634E9, 1.666460682E9, 1.66646073E9, 1.666460778E9, 1.666460826E9, 1.666460874E9, 1.666460922E9, 1.66646097E9, 1.666461018E9, 1.666461066E9, 1.666461114E9, 1.666461162E9, 1.66646121E9, 1.666461258E9, 1.666461306E9, 1.666461354E9, 1.666461402E9, 1.66646145E9, 1.666461498E9, 1.666461546E9, 1.666461594E9, 1.666461642E9, 1.66646169E9, 1.666461738E9, 1.666461786E9, 1.666461834E9, 1.666461882E9, 1.66646193E9, 1.666461978E9, 1.666462026E9, 1.666462074E9, 1.666462122E9, 1.66646217E9, 1.666462218E9, 1.666462266E9, 1.666462314E9, 1.666462362E9, 1.66646241E9, 1.666462458E9, 1.666462506E9, 1.666462554E9, 1.666462602E9, 1.66646265E9, 1.66646304E9, 1.666463041E9, 1.666469028E9, 1.666469076E9, 1.666469124E9, 1.666469172E9, 1.66646922E9, 1.666469268E9, 1.666469316E9, 1.666469364E9, 1.666469412E9, 1.66646946E9, 1.666469508E9, 1.666469556E9, 1.666469604E9, 1.666469652E9, 1.6664697E9, 1.666469748E9, 1.666469796E9, 1.666469844E9, 1.666469892E9, 1.66646994E9, 1.666469988E9, 1.666470036E9, 1.666470084E9, 1.666470132E9, 1.66647018E9, 1.666470228E9, 1.666470276E9, 1.666470324E9, 1.666470372E9, 1.66647042E9, 1.666470468E9, 1.666470516E9, 1.666470564E9, 1.666470612E9, 1.66647066E9, 1.666470708E9, 1.666470756E9, 1.666470804E9, 1.666470852E9, 1.6664709E9, 1.666470948E9, 1.666470996E9, 1.666471044E9, 1.666471092E9, 1.66647114E9, 1.666471188E9, 1.666471236E9, 1.666471284E9, 1.666471332E9, 1.66647138E9, 1.666471428E9, 1.666471476E9, 1.666471524E9, 1.666471572E9, 1.66647162E9, 1.666471668E9, 1.666471716E9, 1.666471764E9, 1.666471812E9, 1.66647186E9, 1.666471908E9, 1.666471956E9, 1.666472004E9, 1.666472052E9, 1.6664721E9, 1.666472148E9, 1.666472196E9, 1.666472244E9, 1.666472292E9, 1.66647234E9, 1.6664727E9, 1.66647288E9, 1.666478707E9, 1.666478755E9, 1.666478803E9, 1.666478851E9, 1.666478899E9, 1.666478947E9, 1.666478995E9, 1.666479043E9, 1.666479091E9, 1.666479139E9, 1.666479187E9, 1.666479235E9, 1.666479283E9, 1.666479331E9, 1.666479379E9, 1.666479427E9, 1.666479475E9, 1.666479523E9, 1.666479571E9, 1.666479619E9, 1.666479667E9, 1.666479715E9, 1.666479763E9, 1.666479811E9, 1.666479859E9, 1.666479907E9, 1.666479955E9, 1.666480003E9, 1.666480051E9, 1.666480099E9, 1.666480147E9, 1.666480195E9, 1.666480243E9, 1.666480291E9, 1.666480339E9, 1.666480387E9, 1.666480435E9, 1.666480483E9, 1.666480531E9, 1.666480579E9, 1.666480627E9, 1.666480675E9, 1.666480723E9, 1.666480771E9, 1.666480819E9, 1.666480867E9, 1.666480915E9, 1.666480963E9, 1.666481011E9, 1.666481059E9, 1.666481107E9, 1.666481155E9, 1.666481203E9, 1.666481251E9, 1.666481299E9, 1.666481347E9, 1.666481395E9, 1.666481443E9, 1.666481491E9, 1.666481539E9, 1.666481587E9, 1.666481635E9, 1.666481683E9, 1.666481731E9, 1.666481779E9, 1.666481827E9, 1.666481875E9, 1.666481923E9, 1.666481971E9, 1.666482019E9, 1.666482067E9, 1.666482115E9, 1.666482163E9, 1.666482211E9, 1.666482259E9, 1.66648254E9, 1.66648272E9, 1.66648845E9, 1.666488498E9, 1.666488546E9, 1.666488594E9, 1.666488642E9, 1.66648869E9, 1.666488738E9, 1.666488786E9, 1.666488834E9, 1.666488882E9, 1.66648893E9, 1.666488978E9, 1.666489026E9, 1.666489074E9, 1.666489122E9, 1.66648917E9, 1.666489218E9, 1.666489266E9, 1.666489314E9, 1.666489362E9, 1.66648941E9, 1.666489458E9, 1.666489506E9, 1.666489554E9, 1.666489602E9, 1.66648965E9, 1.666489698E9, 1.666489746E9, 1.666489794E9, 1.666489842E9, 1.66648989E9, 1.666489938E9, 1.666489986E9, 1.666490034E9, 1.666490082E9, 1.66649013E9, 1.666490178E9, 1.666490226E9, 1.666490274E9, 1.666490322E9, 1.66649037E9, 1.666490418E9, 1.666490466E9, 1.666490514E9, 1.666490562E9, 1.66649061E9, 1.666490658E9, 1.666490706E9, 1.666490754E9, 1.666490802E9, 1.66649085E9, 1.666490898E9, 1.666490946E9, 1.666490994E9, 1.666491042E9, 1.66649109E9, 1.666491138E9, 1.666491186E9, 1.666491234E9, 1.666491282E9, 1.66649133E9, 1.666491378E9, 1.666491426E9, 1.666491474E9, 1.666491522E9, 1.66649157E9, 1.666491618E9, 1.666491666E9, 1.666491714E9, 1.666491762E9, 1.66649181E9, 1.66649214E9, 1.66649232E9, 1.666497916E9, 1.666497964E9, 1.666498012E9, 1.66649806E9, 1.666498108E9, 1.666498156E9, 1.666498204E9, 1.666498252E9, 1.6664983E9, 1.666498348E9, 1.666498396E9, 1.666498444E9, 1.666498492E9, 1.66649854E9, 1.666498588E9, 1.666498636E9, 1.666498684E9, 1.666498732E9, 1.66649878E9, 1.666498828E9, 1.666498876E9, 1.666498924E9, 1.666498972E9, 1.66649902E9, 1.666499068E9, 1.666499116E9, 1.666499164E9, 1.666499212E9, 1.66649926E9, 1.666499308E9, 1.666499356E9, 1.666499404E9, 1.666499452E9, 1.6664995E9, 1.666499548E9, 1.666499596E9, 1.666499644E9, 1.666499692E9, 1.66649974E9, 1.666499788E9, 1.666499836E9, 1.666499884E9, 1.666499932E9, 1.66649998E9, 1.666500028E9, 1.666500076E9, 1.666500124E9, 1.666500172E9, 1.66650022E9, 1.666500268E9, 1.666500316E9, 1.666500364E9, 1.666500412E9, 1.66650046E9, 1.666500508E9, 1.666500556E9, 1.666500604E9, 1.666500652E9, 1.6665007E9, 1.666500748E9, 1.666500796E9, 1.666500844E9, 1.666500892E9, 1.66650094E9, 1.666500988E9, 1.666501036E9, 1.666501084E9, 1.666501132E9, 1.66650118E9, 1.66650156E9, 1.66650174E9, 1.666507832E9, 1.66650788E9, 1.666507928E9, 1.666507976E9, 1.666508024E9, 1.666508072E9, 1.66650812E9, 1.666508168E9, 1.666508216E9, 1.666508264E9, 1.666508312E9, 1.66650836E9, 1.666508408E9, 1.666508456E9, 1.666508504E9, 1.666508552E9, 1.6665086E9, 1.666508648E9, 1.666508696E9, 1.666508744E9, 1.666508792E9, 1.66650884E9, 1.666508888E9, 1.666508936E9, 1.666508984E9, 1.666509032E9, 1.66650908E9, 1.666509128E9, 1.666509176E9, 1.666509224E9, 1.666509272E9, 1.66650932E9, 1.666509368E9, 1.666509416E9, 1.666509464E9, 1.666509512E9, 1.66650956E9, 1.666509608E9, 1.666509656E9, 1.666509704E9, 1.666509752E9, 1.6665098E9, 1.666509848E9, 1.666509896E9, 1.666509944E9, 1.666509992E9, 1.66651004E9, 1.666510088E9, 1.666510136E9, 1.666510184E9, 1.666510232E9, 1.66651028E9, 1.666510328E9, 1.666510376E9, 1.666510424E9, 1.666510472E9, 1.66651052E9, 1.666510568E9, 1.666510616E9, 1.666510664E9, 1.666510712E9, 1.66651076E9, 1.666510808E9, 1.666510856E9, 1.666510904E9, 1.666510952E9, 1.666511E9, 1.666511048E9, 1.666511096E9, 1.666511144E9, 1.666511192E9, 1.66651124E9, 1.66651164E9, 1.666511641E9, 1.666517393E9, 1.666517441E9, 1.666517489E9, 1.666517537E9, 1.666517585E9, 1.666517633E9, 1.666517681E9, 1.666517729E9, 1.666517777E9, 1.666517825E9, 1.666517873E9, 1.666517921E9, 1.666517969E9, 1.666518017E9, 1.666518065E9, 1.666518113E9, 1.666518161E9, 1.666518209E9, 1.666518257E9, 1.666518305E9, 1.666518353E9, 1.666518401E9, 1.666518449E9, 1.666518497E9, 1.666518545E9, 1.666518593E9, 1.666518641E9, 1.666518689E9, 1.666518737E9, 1.666518785E9, 1.666518833E9, 1.666518881E9, 1.666518929E9, 1.666518977E9, 1.666519025E9, 1.666519073E9, 1.666519121E9, 1.666519169E9, 1.666519217E9, 1.666519265E9, 1.666519313E9, 1.666519361E9, 1.666519409E9, 1.666519457E9, 1.666519505E9, 1.666519553E9, 1.666519601E9, 1.666519649E9, 1.666519697E9, 1.666519745E9, 1.666519793E9, 1.666519841E9, 1.666519889E9, 1.666519937E9, 1.666519985E9, 1.666520033E9, 1.666520081E9, 1.666520129E9, 1.666520177E9, 1.666520225E9, 1.666520273E9, 1.666520321E9, 1.666520369E9, 1.666520417E9, 1.666520465E9, 1.666520513E9, 1.666520561E9, 1.666520609E9, 1.666520657E9, 1.666520705E9, 1.666520753E9, 1.666520801E9, 1.666520849E9, 1.66652124E9, 1.66652142E9, 1.666527191E9, 1.666527239E9, 1.666527287E9, 1.666527335E9, 1.666527383E9, 1.666527431E9, 1.666527479E9, 1.666527527E9, 1.666527575E9, 1.666527623E9, 1.666527671E9, 1.666527719E9, 1.666527767E9, 1.666527815E9, 1.666527863E9, 1.666527911E9, 1.666527959E9, 1.666528007E9, 1.666528055E9, 1.666528103E9, 1.666528151E9, 1.666528199E9, 1.666528247E9, 1.666528295E9, 1.666528343E9, 1.666528391E9, 1.666528439E9, 1.666528487E9, 1.666528535E9, 1.666528583E9, 1.666528631E9, 1.666528679E9, 1.666528727E9, 1.666528775E9, 1.666528823E9, 1.666528871E9, 1.666528919E9, 1.666528967E9, 1.666529015E9, 1.666529063E9, 1.666529111E9, 1.666529159E9, 1.666529207E9, 1.666529255E9, 1.666529303E9, 1.666529351E9, 1.666529399E9, 1.666529447E9, 1.666529495E9, 1.666529543E9, 1.666529591E9, 1.666529639E9, 1.666529687E9, 1.666529735E9, 1.666529783E9, 1.666529831E9, 1.666529879E9, 1.666529927E9, 1.666529975E9, 1.666530023E9, 1.666530071E9, 1.666530119E9, 1.666530167E9, 1.666530215E9, 1.666530263E9, 1.666530311E9, 1.666530359E9, 1.666530407E9, 1.666530455E9, 1.666530503E9, 1.666530551E9, 1.666530599E9, 1.66653096E9, 1.66653114E9, 1.666536826E9, 1.666536874E9, 1.666536922E9, 1.66653697E9, 1.666537018E9, 1.666537066E9, 1.666537114E9, 1.666537162E9, 1.66653721E9, 1.666537258E9, 1.666537306E9, 1.666537354E9, 1.666537402E9, 1.66653745E9, 1.666537498E9, 1.666537546E9, 1.666537594E9, 1.666537642E9, 1.66653769E9, 1.666537738E9, 1.666537786E9, 1.666537834E9, 1.666537882E9, 1.66653793E9, 1.666537978E9, 1.666538026E9, 1.666538074E9, 1.666538122E9, 1.66653817E9, 1.666538218E9, 1.666538266E9, 1.666538314E9, 1.666538362E9, 1.66653841E9, 1.666538458E9, 1.666538506E9, 1.666538554E9, 1.666538602E9, 1.66653865E9, 1.666538698E9, 1.666538746E9, 1.666538794E9, 1.666538842E9, 1.66653889E9, 1.666538938E9, 1.666538986E9, 1.666539034E9, 1.666539082E9, 1.66653913E9, 1.666539178E9, 1.666539226E9, 1.666539274E9, 1.666539322E9, 1.66653937E9, 1.666539418E9, 1.666539466E9, 1.666539514E9, 1.666539562E9, 1.66653961E9, 1.666539658E9, 1.666539706E9, 1.666539754E9, 1.666539802E9, 1.66653985E9, 1.666539898E9, 1.666539946E9, 1.666539994E9, 1.666540042E9, 1.66654009E9, 1.66654038E9, 1.66654056E9, 1.666546346E9, 1.666546394E9, 1.666546442E9, 1.66654649E9, 1.666546538E9, 1.666546586E9, 1.666546634E9, 1.666546682E9, 1.66654673E9, 1.666546778E9, 1.666546826E9, 1.666546874E9, 1.666546922E9, 1.66654697E9, 1.666547018E9, 1.666547066E9, 1.666547114E9, 1.666547162E9, 1.66654721E9, 1.666547258E9, 1.666547306E9, 1.666547354E9, 1.666547402E9, 1.66654745E9, 1.666547498E9, 1.666547546E9, 1.666547594E9, 1.666547642E9, 1.66654769E9, 1.666547738E9, 1.666547786E9, 1.666547834E9, 1.666547882E9, 1.66654793E9, 1.666547978E9, 1.666548026E9, 1.666548074E9, 1.666548122E9, 1.66654817E9, 1.666548218E9, 1.666548266E9, 1.666548314E9, 1.666548362E9, 1.66654841E9, 1.666548458E9, 1.666548506E9, 1.666548554E9, 1.666548602E9, 1.66654865E9, 1.666548698E9, 1.666548746E9, 1.666548794E9, 1.666548842E9, 1.66654889E9, 1.666548938E9, 1.666548986E9, 1.666549034E9, 1.666549082E9, 1.66654913E9, 1.666549178E9, 1.666549226E9, 1.666549274E9, 1.666549322E9, 1.66654937E9, 1.666549418E9, 1.666549466E9, 1.666549514E9, 1.666549562E9, 1.66654961E9, 1.66654998E9, 1.66655016E9, 1.666555946E9, 1.666555994E9, 1.666556042E9, 1.66655609E9, 1.666556138E9, 1.666556186E9, 1.666556234E9, 1.666556282E9, 1.66655633E9, 1.666556378E9, 1.666556426E9, 1.666556474E9, 1.666556522E9, 1.66655657E9, 1.666556618E9, 1.666556666E9, 1.666556714E9, 1.666556762E9, 1.66655681E9, 1.666556858E9, 1.666556906E9, 1.666556954E9, 1.666557002E9, 1.66655705E9, 1.666557098E9, 1.666557146E9, 1.666557194E9, 1.666557242E9, 1.66655729E9, 1.666557338E9, 1.666557386E9, 1.666557434E9, 1.666557482E9, 1.66655753E9, 1.666557578E9, 1.666557626E9, 1.666557674E9, 1.666557722E9, 1.66655777E9, 1.666557818E9, 1.666557866E9, 1.666557914E9, 1.666557962E9, 1.66655801E9, 1.666558058E9, 1.666558106E9, 1.666558154E9, 1.666558202E9, 1.66655825E9, 1.666558298E9, 1.666558346E9, 1.666558394E9, 1.666558442E9, 1.66655849E9, 1.666558538E9, 1.666558586E9, 1.666558634E9, 1.666558682E9, 1.66655873E9, 1.666558778E9, 1.666558826E9, 1.666558874E9, 1.666558922E9, 1.66655897E9, 1.666559018E9, 1.666559066E9, 1.666559114E9, 1.666559162E9, 1.66655921E9, 1.666559258E9, 1.666559306E9, 1.666559354E9, 1.666559402E9, 1.66655945E9, 1.66655976E9, 1.66655994E9, 1.666565682E9, 1.66656573E9, 1.666565778E9, 1.666565826E9, 1.666565874E9, 1.666565922E9, 1.66656597E9, 1.666566018E9, 1.666566066E9, 1.666566114E9, 1.666566162E9, 1.66656621E9, 1.666566258E9, 1.666566306E9, 1.666566354E9, 1.666566402E9, 1.66656645E9, 1.666566498E9, 1.666566546E9, 1.666566594E9, 1.666566642E9, 1.66656669E9, 1.666566738E9, 1.666566786E9, 1.666566834E9, 1.666566882E9, 1.66656693E9, 1.666566978E9, 1.666567026E9, 1.666567074E9, 1.666567122E9, 1.66656717E9, 1.666567218E9, 1.666567266E9, 1.666567314E9, 1.666567362E9, 1.66656741E9, 1.666567458E9, 1.666567506E9, 1.666567554E9, 1.666567602E9, 1.66656765E9, 1.666567698E9, 1.666567746E9, 1.666567794E9, 1.666567842E9, 1.66656789E9, 1.666567938E9, 1.666567986E9, 1.666568034E9, 1.666568082E9, 1.66656813E9, 1.666568178E9, 1.666568226E9, 1.666568274E9, 1.666568322E9, 1.66656837E9, 1.666568418E9, 1.666568466E9, 1.666568514E9, 1.666568562E9, 1.66656861E9, 1.666568658E9, 1.666568706E9, 1.666568754E9, 1.666568802E9, 1.66656885E9, 1.666568898E9, 1.666568946E9, 1.666568994E9, 1.666569042E9, 1.66656909E9, 1.66656936E9, 1.666569361E9, 1.666575247E9, 1.666575295E9, 1.666575343E9, 1.666575391E9, 1.666575439E9, 1.666575487E9, 1.666575535E9, 1.666575583E9, 1.666575631E9, 1.666575679E9, 1.666575727E9, 1.666575775E9, 1.666575823E9, 1.666575871E9, 1.666575919E9, 1.666575967E9, 1.666576015E9, 1.666576063E9, 1.666576111E9, 1.666576159E9, 1.666576207E9, 1.666576255E9, 1.666576303E9, 1.666576351E9, 1.666576399E9, 1.666576447E9, 1.666576495E9, 1.666576543E9, 1.666576591E9, 1.666576639E9, 1.666576687E9, 1.666576735E9, 1.666576783E9, 1.666576831E9, 1.666576879E9, 1.666576927E9, 1.666576975E9, 1.666577023E9, 1.666577071E9, 1.666577119E9, 1.666577167E9, 1.666577215E9, 1.666577263E9, 1.666577311E9, 1.666577359E9, 1.666577407E9, 1.666577455E9, 1.666577503E9, 1.666577551E9, 1.666577599E9, 1.666577647E9, 1.666577695E9, 1.666577743E9, 1.666577791E9, 1.666577839E9, 1.666577887E9, 1.666577935E9, 1.666577983E9, 1.666578031E9, 1.666578079E9, 1.666578127E9, 1.666578175E9, 1.666578223E9, 1.666578271E9, 1.666578319E9, 1.666578367E9, 1.666578415E9, 1.666578463E9, 1.666578511E9, 1.666578559E9, 1.66657896E9, 1.66657926E9, 1.666585052E9, 1.6665851E9, 1.666585148E9, 1.666585196E9, 1.666585244E9, 1.666585292E9, 1.66658534E9, 1.666585388E9, 1.666585436E9, 1.666585484E9, 1.666585532E9, 1.66658558E9, 1.666585628E9, 1.666585676E9, 1.666585724E9, 1.666585772E9, 1.66658582E9, 1.666585868E9, 1.666585916E9, 1.666585964E9, 1.666586012E9, 1.66658606E9, 1.666586108E9, 1.666586156E9, 1.666586204E9, 1.666586252E9, 1.6665863E9, 1.666586348E9, 1.666586396E9, 1.666586444E9, 1.666586492E9, 1.66658654E9, 1.666586588E9, 1.666586636E9, 1.666586684E9, 1.666586732E9, 1.66658678E9, 1.666586828E9, 1.666586876E9, 1.666586924E9, 1.666586972E9, 1.66658702E9, 1.666587068E9, 1.666587116E9, 1.666587164E9, 1.666587212E9, 1.66658726E9, 1.666587308E9, 1.666587356E9, 1.666587404E9, 1.666587452E9, 1.6665875E9, 1.666587548E9, 1.666587596E9, 1.666587644E9, 1.666587692E9, 1.66658774E9, 1.666587788E9, 1.666587836E9, 1.666587884E9, 1.666587932E9, 1.66658798E9, 1.666588028E9, 1.666588076E9, 1.666588124E9, 1.666588172E9, 1.66658822E9, 1.666588268E9, 1.666588316E9, 1.666588364E9, 1.666588412E9, 1.66658846E9, 1.6665888E9, 1.66658904E9, 1.666594679E9, 1.666594727E9, 1.666594775E9, 1.666594823E9, 1.666594871E9, 1.666594919E9, 1.666594967E9, 1.666595015E9, 1.666595063E9, 1.666595111E9, 1.666595159E9, 1.666595207E9, 1.666595255E9, 1.666595303E9, 1.666595351E9, 1.666595399E9, 1.666595447E9, 1.666595495E9, 1.666595543E9, 1.666595591E9, 1.666595639E9, 1.666595687E9, 1.666595735E9, 1.666595783E9, 1.666595831E9, 1.666595879E9, 1.666595927E9, 1.666595975E9, 1.666596023E9, 1.666596071E9, 1.666596119E9, 1.666596167E9, 1.666596215E9, 1.666596263E9, 1.666596311E9, 1.666596359E9, 1.666596407E9, 1.666596455E9, 1.666596503E9, 1.666596551E9, 1.666596599E9, 1.666596647E9, 1.666596695E9, 1.666596743E9, 1.666596791E9, 1.666596839E9, 1.666596887E9, 1.666596935E9, 1.666596983E9, 1.666597031E9, 1.666597079E9, 1.666597127E9, 1.666597175E9, 1.666597223E9, 1.666597271E9, 1.666597319E9, 1.666597367E9, 1.666597415E9, 1.666597463E9, 1.666597511E9, 1.666597559E9, 1.666597607E9, 1.666597655E9, 1.666597703E9, 1.666597751E9, 1.666597799E9, 1.666597847E9, 1.666597895E9, 1.666597943E9, 1.666597991E9, 1.666598039E9, 1.66659846E9, 1.66659864E9, 1.666604539E9, 1.666604587E9, 1.666604635E9, 1.666604683E9, 1.666604731E9, 1.666604779E9, 1.666604827E9, 1.666604875E9, 1.666604923E9, 1.666604971E9, 1.666605019E9, 1.666605067E9, 1.666605115E9, 1.666605163E9, 1.666605211E9, 1.666605259E9, 1.666605307E9, 1.666605355E9, 1.666605403E9, 1.666605451E9, 1.666605499E9, 1.666605547E9, 1.666605595E9, 1.666605643E9, 1.666605691E9, 1.666605739E9, 1.666605787E9, 1.666605835E9, 1.666605883E9, 1.666605931E9, 1.666605979E9, 1.666606027E9, 1.666606075E9, 1.666606123E9, 1.666606171E9, 1.666606219E9, 1.666606267E9, 1.666606315E9, 1.666606363E9, 1.666606411E9, 1.666606459E9, 1.666606507E9, 1.666606555E9, 1.666606603E9, 1.666606651E9, 1.666606699E9, 1.666606747E9, 1.666606795E9, 1.666606843E9, 1.666606891E9, 1.666606939E9, 1.666606987E9, 1.666607035E9, 1.666607083E9, 1.666607131E9, 1.666607179E9, 1.666607227E9, 1.666607275E9, 1.666607323E9, 1.666607371E9, 1.666607419E9, 1.666607467E9, 1.666607515E9, 1.666607563E9, 1.666607611E9, 1.666607659E9, 1.666607707E9, 1.666607755E9, 1.666607803E9, 1.666607851E9, 1.666607899E9, 1.6666083E9, 1.66660848E9, 1.666614197E9, 1.666614245E9, 1.666614293E9, 1.666614341E9, 1.666614389E9, 1.666614437E9, 1.666614485E9, 1.666614533E9, 1.666614581E9, 1.666614629E9, 1.666614677E9, 1.666614725E9, 1.666614773E9, 1.666614821E9, 1.666614869E9, 1.666614917E9, 1.666614965E9, 1.666615013E9, 1.666615061E9, 1.666615109E9, 1.666615157E9, 1.666615205E9, 1.666615253E9, 1.666615301E9, 1.666615349E9, 1.666615397E9, 1.666615445E9, 1.666615493E9, 1.666615541E9, 1.666615589E9, 1.666615637E9, 1.666615685E9, 1.666615733E9, 1.666615781E9, 1.666615829E9, 1.666615877E9, 1.666615925E9, 1.666615973E9, 1.666616021E9, 1.666616069E9, 1.666616117E9, 1.666616165E9, 1.666616213E9, 1.666616261E9, 1.666616309E9, 1.666616357E9, 1.666616405E9, 1.666616453E9, 1.666616501E9, 1.666616549E9, 1.666616597E9, 1.666616645E9, 1.666616693E9, 1.666616741E9, 1.666616789E9, 1.666616837E9, 1.666616885E9, 1.666616933E9, 1.666616981E9, 1.666617029E9, 1.666617077E9, 1.666617125E9, 1.666617173E9, 1.666617221E9, 1.666617269E9, 1.666617317E9, 1.666617365E9, 1.666617413E9, 1.666617461E9, 1.666617509E9, 1.6666179E9, 1.66661808E9, 1.666623912E9, 1.66662396E9, 1.666624008E9, 1.666624056E9, 1.666624104E9, 1.666624152E9, 1.6666242E9, 1.666624248E9, 1.666624296E9, 1.666624344E9, 1.666624392E9, 1.66662444E9, 1.666624488E9, 1.666624536E9, 1.666624584E9, 1.666624632E9, 1.66662468E9, 1.666624728E9, 1.666624776E9, 1.666624824E9, 1.666624872E9, 1.66662492E9, 1.666624968E9, 1.666625016E9, 1.666625064E9, 1.666625112E9, 1.66662516E9, 1.666625208E9, 1.666625256E9, 1.666625304E9, 1.666625352E9, 1.6666254E9, 1.666625448E9, 1.666625496E9, 1.666625544E9, 1.666625592E9, 1.66662564E9, 1.666625688E9, 1.666625736E9, 1.666625784E9, 1.666625832E9, 1.66662588E9, 1.666625928E9, 1.666625976E9, 1.666626024E9, 1.666626072E9, 1.66662612E9, 1.666626168E9, 1.666626216E9, 1.666626264E9, 1.666626312E9, 1.66662636E9, 1.666626408E9, 1.666626456E9, 1.666626504E9, 1.666626552E9, 1.6666266E9, 1.666626648E9, 1.666626696E9, 1.666626744E9, 1.666626792E9, 1.66662684E9, 1.666626888E9, 1.666626936E9, 1.666626984E9, 1.666627032E9, 1.66662708E9, 1.666627128E9, 1.666627176E9, 1.666627224E9, 1.666627272E9, 1.66662732E9, 1.66662762E9, 1.6666278E9, 1.666633534E9, 1.666633582E9, 1.66663363E9, 1.666633678E9, 1.666633726E9, 1.666633774E9, 1.666633822E9, 1.66663387E9, 1.666633918E9, 1.666633966E9, 1.666634014E9, 1.666634062E9, 1.66663411E9, 1.666634158E9, 1.666634206E9, 1.666634254E9, 1.666634302E9, 1.66663435E9, 1.666634398E9, 1.666634446E9, 1.666634494E9, 1.666634542E9, 1.66663459E9, 1.666634638E9, 1.666634686E9, 1.666634734E9, 1.666634782E9, 1.66663483E9, 1.666634878E9, 1.666634926E9, 1.666634974E9, 1.666635022E9, 1.66663507E9, 1.666635118E9, 1.666635166E9, 1.666635214E9, 1.666635262E9, 1.66663531E9, 1.666635358E9, 1.666635406E9, 1.666635454E9, 1.666635502E9, 1.66663555E9, 1.666635598E9, 1.666635646E9, 1.666635694E9, 1.666635742E9, 1.66663579E9, 1.666635838E9, 1.666635886E9, 1.666635934E9, 1.666635982E9, 1.66663603E9, 1.666636078E9, 1.666636126E9, 1.666636174E9, 1.666636222E9, 1.66663627E9, 1.666636318E9, 1.666636366E9, 1.666636414E9, 1.666636462E9, 1.66663651E9, 1.666636558E9, 1.666636606E9, 1.666636654E9, 1.666636702E9, 1.66663675E9, 1.66663704E9, 1.66663722E9, 1.666642952E9, 1.666643E9, 1.666643048E9, 1.666643096E9, 1.666643144E9, 1.666643192E9, 1.66664324E9, 1.666643288E9, 1.666643336E9, 1.666643384E9, 1.666643432E9, 1.66664348E9, 1.666643528E9, 1.666643576E9, 1.666643624E9, 1.666643672E9, 1.66664372E9, 1.666643768E9, 1.666643816E9, 1.666643864E9, 1.666643912E9, 1.66664396E9, 1.666644008E9, 1.666644056E9, 1.666644104E9, 1.666644152E9, 1.6666442E9, 1.666644248E9, 1.666644296E9, 1.666644344E9, 1.666644392E9, 1.66664444E9, 1.666644488E9, 1.666644536E9, 1.666644584E9, 1.666644632E9, 1.66664468E9, 1.666644728E9, 1.666644776E9, 1.666644824E9, 1.666644872E9, 1.66664492E9, 1.666644968E9, 1.666645016E9, 1.666645064E9, 1.666645112E9, 1.66664516E9, 1.666645208E9, 1.666645256E9, 1.666645304E9, 1.666645352E9, 1.6666454E9, 1.666645448E9, 1.666645496E9, 1.666645544E9, 1.666645592E9, 1.66664564E9, 1.666645688E9, 1.666645736E9, 1.666645784E9, 1.666645832E9, 1.66664588E9, 1.666645928E9, 1.666645976E9, 1.666646024E9, 1.666646072E9, 1.66664612E9, 1.666646168E9, 1.666646216E9, 1.666646264E9, 1.666646312E9, 1.66664636E9, 1.66664664E9, 1.66664682E9, 1.666652635E9, 1.666652683E9, 1.666652731E9, 1.666652779E9, 1.666652827E9, 1.666652875E9, 1.666652923E9, 1.666652971E9, 1.666653019E9, 1.666653067E9, 1.666653115E9, 1.666653163E9, 1.666653211E9, 1.666653259E9, 1.666653307E9, 1.666653355E9, 1.666653403E9, 1.666653451E9, 1.666653499E9, 1.666653547E9, 1.666653595E9, 1.666653643E9, 1.666653691E9, 1.666653739E9, 1.666653787E9, 1.666653835E9, 1.666653883E9, 1.666653931E9, 1.666653979E9, 1.666654027E9, 1.666654075E9, 1.666654123E9, 1.666654171E9, 1.666654219E9, 1.666654267E9, 1.666654315E9, 1.666654363E9, 1.666654411E9, 1.666654459E9, 1.666654507E9, 1.666654555E9, 1.666654603E9, 1.666654651E9, 1.666654699E9, 1.666654747E9, 1.666654795E9, 1.666654843E9, 1.666654891E9, 1.666654939E9, 1.666654987E9, 1.666655035E9, 1.666655083E9, 1.666655131E9, 1.666655179E9, 1.666655227E9, 1.666655275E9, 1.666655323E9, 1.666655371E9, 1.666655419E9, 1.666655467E9, 1.666655515E9, 1.666655563E9, 1.666655611E9, 1.666655659E9, 1.666655707E9, 1.666655755E9, 1.666655803E9, 1.666655851E9, 1.666655899E9, 1.66665624E9, 1.66665642E9, 1.666662443E9, 1.666662491E9, 1.666662539E9, 1.666662587E9, 1.666662635E9, 1.666662683E9, 1.666662731E9, 1.666662779E9, 1.666662827E9, 1.666662875E9, 1.666662923E9, 1.666662971E9, 1.666663019E9, 1.666663067E9, 1.666663115E9, 1.666663163E9, 1.666663211E9, 1.666663259E9, 1.666663307E9, 1.666663355E9, 1.666663403E9, 1.666663451E9, 1.666663499E9, 1.666663547E9, 1.666663595E9, 1.666663643E9, 1.666663691E9, 1.666663739E9, 1.666663787E9, 1.666663835E9, 1.666663883E9, 1.666663931E9, 1.666663979E9, 1.666664027E9, 1.666664075E9, 1.666664123E9, 1.666664171E9, 1.666664219E9, 1.666664267E9, 1.666664315E9, 1.666664363E9, 1.666664411E9, 1.666664459E9, 1.666664507E9, 1.666664555E9, 1.666664603E9, 1.666664651E9, 1.666664699E9, 1.666664747E9, 1.666664795E9, 1.666664843E9, 1.666664891E9, 1.666664939E9, 1.666664987E9, 1.666665035E9, 1.666665083E9, 1.666665131E9, 1.666665179E9, 1.666665227E9, 1.666665275E9, 1.666665323E9, 1.666665371E9, 1.666665419E9, 1.666665467E9, 1.666665515E9, 1.666665563E9, 1.666665611E9, 1.666665659E9, 1.666665707E9, 1.666665755E9, 1.666665803E9, 1.666665851E9, 1.666665899E9, 1.6666662E9, 1.66666638E9, 1.666672181E9, 1.666672229E9, 1.666672277E9, 1.666672325E9, 1.666672373E9, 1.666672421E9, 1.666672469E9, 1.666672517E9, 1.666672565E9, 1.666672613E9, 1.666672661E9, 1.666672709E9, 1.666672757E9, 1.666672805E9, 1.666672853E9, 1.666672901E9, 1.666672949E9, 1.666672997E9, 1.666673045E9, 1.666673093E9, 1.666673141E9, 1.666673189E9, 1.666673237E9, 1.666673285E9, 1.666673333E9, 1.666673381E9, 1.666673429E9, 1.666673477E9, 1.666673525E9, 1.666673573E9, 1.666673621E9, 1.666673669E9, 1.666673717E9, 1.666673765E9, 1.666673813E9, 1.666673861E9, 1.666673909E9, 1.666673957E9, 1.666674005E9, 1.666674053E9, 1.666674101E9, 1.666674149E9, 1.666674197E9, 1.666674245E9, 1.666674293E9, 1.666674341E9, 1.666674389E9, 1.666674437E9, 1.666674485E9, 1.666674533E9, 1.666674581E9, 1.666674629E9, 1.666674677E9, 1.666674725E9, 1.666674773E9, 1.666674821E9, 1.666674869E9, 1.666674917E9, 1.666674965E9, 1.666675013E9, 1.666675061E9, 1.666675109E9, 1.666675157E9, 1.666675205E9, 1.666675253E9, 1.666675301E9, 1.666675349E9, 1.666675397E9, 1.666675445E9, 1.666675493E9, 1.666675541E9, 1.666675589E9, 1.66667592E9, 1.6666761E9, 1.666681863E9, 1.666681911E9, 1.666681959E9, 1.666682007E9, 1.666682055E9, 1.666682103E9, 1.666682151E9, 1.666682199E9, 1.666682247E9, 1.666682295E9, 1.666682343E9, 1.666682391E9, 1.666682439E9, 1.666682487E9, 1.666682535E9, 1.666682583E9, 1.666682631E9, 1.666682679E9, 1.666682727E9, 1.666682775E9, 1.666682823E9, 1.666682871E9, 1.666682919E9, 1.666682967E9, 1.666683015E9, 1.666683063E9, 1.666683111E9, 1.666683159E9, 1.666683207E9, 1.666683255E9, 1.666683303E9, 1.666683351E9, 1.666683399E9, 1.666683447E9, 1.666683495E9, 1.666683543E9, 1.666683591E9, 1.666683639E9, 1.666683687E9, 1.666683735E9, 1.666683783E9, 1.666683831E9, 1.666683879E9, 1.666683927E9, 1.666683975E9, 1.666684023E9, 1.666684071E9, 1.666684119E9, 1.666684167E9, 1.666684215E9, 1.666684263E9, 1.666684311E9, 1.666684359E9, 1.666684407E9, 1.666684455E9, 1.666684503E9, 1.666684551E9, 1.666684599E9, 1.666684647E9, 1.666684695E9, 1.666684743E9, 1.666684791E9, 1.666684839E9, 1.666684887E9, 1.666684935E9, 1.666684983E9, 1.666685031E9, 1.666685079E9, 1.6666854E9, 1.66668558E9, 1.66669121E9, 1.666691258E9, 1.666691306E9, 1.666691354E9, 1.666691402E9, 1.66669145E9, 1.666691498E9, 1.666691546E9, 1.666691594E9, 1.666691642E9, 1.66669169E9, 1.666691738E9, 1.666691786E9, 1.666691834E9, 1.666691882E9, 1.66669193E9, 1.666691978E9, 1.666692026E9, 1.666692074E9, 1.666692122E9, 1.66669217E9, 1.666692218E9, 1.666692266E9, 1.666692314E9, 1.666692362E9, 1.66669241E9, 1.666692458E9, 1.666692506E9, 1.666692554E9, 1.666692602E9, 1.66669265E9, 1.666692698E9, 1.666692746E9, 1.666692794E9, 1.666692842E9, 1.66669289E9, 1.666692938E9, 1.666692986E9, 1.666693034E9, 1.666693082E9, 1.66669313E9, 1.666693178E9, 1.666693226E9, 1.666693274E9, 1.666693322E9, 1.66669337E9, 1.666693418E9, 1.666693466E9, 1.666693514E9, 1.666693562E9, 1.66669361E9, 1.666693658E9, 1.666693706E9, 1.666693754E9, 1.666693802E9, 1.66669385E9, 1.666693898E9, 1.666693946E9, 1.666693994E9, 1.666694042E9, 1.66669409E9, 1.666694138E9, 1.666694186E9, 1.666694234E9, 1.666694282E9, 1.66669433E9, 1.666694378E9, 1.666694426E9, 1.666694474E9, 1.666694522E9, 1.66669457E9, 1.66669494E9, 1.66669512E9, 1.666700818E9, 1.666700866E9, 1.666700914E9, 1.666700962E9, 1.66670101E9, 1.666701058E9, 1.666701106E9, 1.666701154E9, 1.666701202E9, 1.66670125E9, 1.666701298E9, 1.666701346E9, 1.666701394E9, 1.666701442E9, 1.66670149E9, 1.666701538E9, 1.666701586E9, 1.666701634E9, 1.666701682E9, 1.66670173E9, 1.666701778E9, 1.666701826E9, 1.666701874E9, 1.666701922E9, 1.66670197E9, 1.666702018E9, 1.666702066E9, 1.666702114E9, 1.666702162E9, 1.66670221E9, 1.666702258E9, 1.666702306E9, 1.666702354E9, 1.666702402E9, 1.66670245E9, 1.666702498E9, 1.666702546E9, 1.666702594E9, 1.666702642E9, 1.66670269E9, 1.666702738E9, 1.666702786E9, 1.666702834E9, 1.666702882E9, 1.66670293E9, 1.666702978E9, 1.666703026E9, 1.666703074E9, 1.666703122E9, 1.66670317E9, 1.666703218E9, 1.666703266E9, 1.666703314E9, 1.666703362E9, 1.66670341E9, 1.666703458E9, 1.666703506E9, 1.666703554E9, 1.666703602E9, 1.66670365E9, 1.666703698E9, 1.666703746E9, 1.666703794E9, 1.666703842E9, 1.66670389E9, 1.666703938E9, 1.666703986E9, 1.666704034E9, 1.666704082E9, 1.66670413E9, 1.66670442E9, 1.6667046E9, 1.66671034E9, 1.666710388E9, 1.666710436E9, 1.666710484E9, 1.666710532E9, 1.66671058E9, 1.666710628E9, 1.666710676E9, 1.666710724E9, 1.666710772E9, 1.66671082E9, 1.666710868E9, 1.666710916E9, 1.666710964E9, 1.666711012E9, 1.66671106E9, 1.666711108E9, 1.666711156E9, 1.666711204E9, 1.666711252E9, 1.6667113E9, 1.666711348E9, 1.666711396E9, 1.666711444E9, 1.666711492E9, 1.66671154E9, 1.666711588E9, 1.666711636E9, 1.666711684E9, 1.666711732E9, 1.66671178E9, 1.666711828E9, 1.666711876E9, 1.666711924E9, 1.666711972E9, 1.66671202E9, 1.666712068E9, 1.666712116E9, 1.666712164E9, 1.666712212E9, 1.66671226E9, 1.666712308E9, 1.666712356E9, 1.666712404E9, 1.666712452E9, 1.6667125E9, 1.666712548E9, 1.666712596E9, 1.666712644E9, 1.666712692E9, 1.66671274E9, 1.666712788E9, 1.666712836E9, 1.666712884E9, 1.666712932E9, 1.66671298E9, 1.666713028E9, 1.666713076E9, 1.666713124E9, 1.666713172E9, 1.66671322E9, 1.666713268E9, 1.666713316E9, 1.666713364E9, 1.666713412E9, 1.66671346E9, 1.666713508E9, 1.666713556E9, 1.666713604E9, 1.666713652E9, 1.6667137E9, 1.66671402E9, 1.6667142E9, 1.666719945E9, 1.666719993E9, 1.666720041E9, 1.666720089E9, 1.666720137E9, 1.666720185E9, 1.666720233E9, 1.666720281E9, 1.666720329E9, 1.666720377E9, 1.666720425E9, 1.666720473E9, 1.666720521E9, 1.666720569E9, 1.666720617E9, 1.666720665E9, 1.666720713E9, 1.666720761E9, 1.666720809E9, 1.666720857E9, 1.666720905E9, 1.666720953E9, 1.666721001E9, 1.666721049E9, 1.666721097E9, 1.666721145E9, 1.666721193E9, 1.666721241E9, 1.666721289E9, 1.666721337E9, 1.666721385E9, 1.666721433E9, 1.666721481E9, 1.666721529E9, 1.666721577E9, 1.666721625E9, 1.666721673E9, 1.666721721E9, 1.666721769E9, 1.666721817E9, 1.666721865E9, 1.666721913E9, 1.666721961E9, 1.666722009E9, 1.666722057E9, 1.666722105E9, 1.666722153E9, 1.666722201E9, 1.666722249E9, 1.666722297E9, 1.666722345E9, 1.666722393E9, 1.666722441E9, 1.666722489E9, 1.666722537E9, 1.666722585E9, 1.666722633E9, 1.666722681E9, 1.666722729E9, 1.666722777E9, 1.666722825E9, 1.666722873E9, 1.666722921E9, 1.666722969E9, 1.666723017E9, 1.666723065E9, 1.666723113E9, 1.666723161E9, 1.666723209E9, 1.66672356E9, 1.66672374E9, 1.66672947E9, 1.666729518E9, 1.666729566E9, 1.666729614E9, 1.666729662E9, 1.66672971E9, 1.666729758E9, 1.666729806E9, 1.666729854E9, 1.666729902E9, 1.66672995E9, 1.666729998E9, 1.666730046E9, 1.666730094E9, 1.666730142E9, 1.66673019E9, 1.666730238E9, 1.666730286E9, 1.666730334E9, 1.666730382E9, 1.66673043E9, 1.666730478E9, 1.666730526E9, 1.666730574E9, 1.666730622E9, 1.66673067E9, 1.666730718E9, 1.666730766E9, 1.666730814E9, 1.666730862E9, 1.66673091E9, 1.666730958E9, 1.666731006E9, 1.666731054E9, 1.666731102E9, 1.66673115E9, 1.666731198E9, 1.666731246E9, 1.666731294E9, 1.666731342E9, 1.66673139E9, 1.666731438E9, 1.666731486E9, 1.666731534E9, 1.666731582E9, 1.66673163E9, 1.666731678E9, 1.666731726E9, 1.666731774E9, 1.666731822E9, 1.66673187E9, 1.666731918E9, 1.666731966E9, 1.666732014E9, 1.666732062E9, 1.66673211E9, 1.666732158E9, 1.666732206E9, 1.666732254E9, 1.666732302E9, 1.66673235E9, 1.666732398E9, 1.666732446E9, 1.666732494E9, 1.666732542E9, 1.66673259E9, 1.666732638E9, 1.666732686E9, 1.666732734E9, 1.666732782E9, 1.66673283E9, 1.6667331E9, 1.66673328E9, 1.666738915E9, 1.666738963E9, 1.666739011E9, 1.666739059E9, 1.666739107E9, 1.666739155E9, 1.666739203E9, 1.666739251E9, 1.666739299E9, 1.666739347E9, 1.666739395E9, 1.666739443E9, 1.666739491E9, 1.666739539E9, 1.666739587E9, 1.666739635E9, 1.666739683E9, 1.666739731E9, 1.666739779E9, 1.666739827E9, 1.666739875E9, 1.666739923E9, 1.666739971E9, 1.666740019E9, 1.666740067E9, 1.666740115E9, 1.666740163E9, 1.666740211E9, 1.666740259E9, 1.666740307E9, 1.666740355E9, 1.666740403E9, 1.666740451E9, 1.666740499E9, 1.666740547E9, 1.666740595E9, 1.666740643E9, 1.666740691E9, 1.666740739E9, 1.666740787E9, 1.666740835E9, 1.666740883E9, 1.666740931E9, 1.666740979E9, 1.666741027E9, 1.666741075E9, 1.666741123E9, 1.666741171E9, 1.666741219E9, 1.666741267E9, 1.666741315E9, 1.666741363E9, 1.666741411E9, 1.666741459E9, 1.666741507E9, 1.666741555E9, 1.666741603E9, 1.666741651E9, 1.666741699E9, 1.666741747E9, 1.666741795E9, 1.666741843E9, 1.666741891E9, 1.666741939E9, 1.666741987E9, 1.666742035E9, 1.666742083E9, 1.666742131E9, 1.666742179E9, 1.666742227E9, 1.666742275E9, 1.666742323E9, 1.666742371E9, 1.666742419E9, 1.66674282E9, 1.666743E9, 1.666748883E9, 1.666748931E9, 1.666748979E9, 1.666749027E9, 1.666749075E9, 1.666749123E9, 1.666749171E9, 1.666749219E9, 1.666749267E9, 1.666749315E9, 1.666749363E9, 1.666749411E9, 1.666749459E9, 1.666749507E9, 1.666749555E9, 1.666749603E9, 1.666749651E9, 1.666749699E9, 1.666749747E9, 1.666749795E9, 1.666749843E9, 1.666749891E9, 1.666749939E9, 1.666749987E9, 1.666750035E9, 1.666750083E9, 1.666750131E9, 1.666750179E9, 1.666750227E9, 1.666750275E9, 1.666750323E9, 1.666750371E9, 1.666750419E9, 1.666750467E9, 1.666750515E9, 1.666750563E9, 1.666750611E9, 1.666750659E9, 1.666750707E9, 1.666750755E9, 1.666750803E9, 1.666750851E9, 1.666750899E9, 1.666750947E9, 1.666750995E9, 1.666751043E9, 1.666751091E9, 1.666751139E9, 1.666751187E9, 1.666751235E9, 1.666751283E9, 1.666751331E9, 1.666751379E9, 1.666751427E9, 1.666751475E9, 1.666751523E9, 1.666751571E9, 1.666751619E9, 1.666751667E9, 1.666751715E9, 1.666751763E9, 1.666751811E9, 1.666751859E9, 1.666751907E9, 1.666751955E9, 1.666752003E9, 1.666752051E9, 1.666752099E9, 1.66675242E9, 1.6667526E9, 1.666758229E9, 1.666758277E9, 1.666758325E9, 1.666758373E9, 1.666758421E9, 1.666758469E9, 1.666758517E9, 1.666758565E9, 1.666758613E9, 1.666758661E9, 1.666758709E9, 1.666758757E9, 1.666758805E9, 1.666758853E9, 1.666758901E9, 1.666758949E9, 1.666758997E9, 1.666759045E9, 1.666759093E9, 1.666759141E9, 1.666759189E9, 1.666759237E9, 1.666759285E9, 1.666759333E9, 1.666759381E9, 1.666759429E9, 1.666759477E9, 1.666759525E9, 1.666759573E9, 1.666759621E9, 1.666759669E9, 1.666759717E9, 1.666759765E9, 1.666759813E9, 1.666759861E9, 1.666759909E9, 1.666759957E9, 1.666760005E9, 1.666760053E9, 1.666760101E9, 1.666760149E9, 1.666760197E9, 1.666760245E9, 1.666760293E9, 1.666760341E9, 1.666760389E9, 1.666760437E9, 1.666760485E9, 1.666760533E9, 1.666760581E9, 1.666760629E9, 1.666760677E9, 1.666760725E9, 1.666760773E9, 1.666760821E9, 1.666760869E9, 1.666760917E9, 1.666760965E9, 1.666761013E9, 1.666761061E9, 1.666761109E9, 1.666761157E9, 1.666761205E9, 1.666761253E9, 1.666761301E9, 1.666761349E9, 1.66676166E9, 1.66676184E9, 1.66676768E9, 1.666767728E9, 1.666767776E9, 1.666767824E9, 1.666767872E9, 1.66676792E9, 1.666767968E9, 1.666768016E9, 1.666768064E9, 1.666768112E9, 1.66676816E9, 1.666768208E9, 1.666768256E9, 1.666768304E9, 1.666768352E9, 1.6667684E9, 1.666768448E9, 1.666768496E9, 1.666768544E9, 1.666768592E9, 1.66676864E9, 1.666768688E9, 1.666768736E9, 1.666768784E9, 1.666768832E9, 1.66676888E9, 1.666768928E9, 1.666768976E9, 1.666769024E9, 1.666769072E9, 1.66676912E9, 1.666769168E9, 1.666769216E9, 1.666769264E9, 1.666769312E9, 1.66676936E9, 1.666769408E9, 1.666769456E9, 1.666769504E9, 1.666769552E9, 1.6667696E9, 1.666769648E9, 1.666769696E9, 1.666769744E9, 1.666769792E9, 1.66676984E9, 1.666769888E9, 1.666769936E9, 1.666769984E9, 1.666770032E9, 1.66677008E9, 1.666770128E9, 1.666770176E9, 1.666770224E9, 1.666770272E9, 1.66677032E9, 1.666770368E9, 1.666770416E9, 1.666770464E9, 1.666770512E9, 1.66677056E9, 1.666770608E9, 1.666770656E9, 1.666770704E9, 1.666770752E9, 1.6667708E9, 1.666770848E9, 1.666770896E9, 1.666770944E9, 1.666770992E9, 1.66677104E9, 1.66677138E9, 1.66677156E9, 1.666777423E9, 1.666777471E9, 1.666777519E9, 1.666777567E9, 1.666777615E9, 1.666777663E9, 1.666777711E9, 1.666777759E9, 1.666777807E9, 1.666777855E9, 1.666777903E9, 1.666777951E9, 1.666777999E9, 1.666778047E9, 1.666778095E9, 1.666778143E9, 1.666778191E9, 1.666778239E9, 1.666778287E9, 1.666778335E9, 1.666778383E9, 1.666778431E9, 1.666778479E9, 1.666778527E9, 1.666778575E9, 1.666778623E9, 1.666778671E9, 1.666778719E9, 1.666778767E9, 1.666778815E9, 1.666778863E9, 1.666778911E9, 1.666778959E9, 1.666779007E9, 1.666779055E9, 1.666779103E9, 1.666779151E9, 1.666779199E9, 1.666779247E9, 1.666779295E9, 1.666779343E9, 1.666779391E9, 1.666779439E9, 1.666779487E9, 1.666779535E9, 1.666779583E9, 1.666779631E9, 1.666779679E9, 1.666779727E9, 1.666779775E9, 1.666779823E9, 1.666779871E9, 1.666779919E9, 1.666779967E9, 1.666780015E9, 1.666780063E9, 1.666780111E9, 1.666780159E9, 1.666780207E9, 1.666780255E9, 1.666780303E9, 1.666780351E9, 1.666780399E9, 1.666780447E9, 1.666780495E9, 1.666780543E9, 1.666780591E9, 1.666780639E9, 1.666780687E9, 1.666780735E9, 1.666780783E9, 1.666780831E9, 1.666780879E9, 1.66678122E9, 1.6667814E9, 1.666787138E9, 1.666787186E9, 1.666787234E9, 1.666787282E9, 1.66678733E9, 1.666787378E9, 1.666787426E9, 1.666787474E9, 1.666787522E9, 1.66678757E9, 1.666787618E9, 1.666787666E9, 1.666787714E9, 1.666787762E9, 1.66678781E9, 1.666787858E9, 1.666787906E9, 1.666787954E9, 1.666788002E9, 1.66678805E9, 1.666788098E9, 1.666788146E9, 1.666788194E9, 1.666788242E9, 1.66678829E9, 1.666788338E9, 1.666788386E9, 1.666788434E9, 1.666788482E9, 1.66678853E9, 1.666788578E9, 1.666788626E9, 1.666788674E9, 1.666788722E9, 1.66678877E9, 1.666788818E9, 1.666788866E9, 1.666788914E9, 1.666788962E9, 1.66678901E9, 1.666789058E9, 1.666789106E9, 1.666789154E9, 1.666789202E9, 1.66678925E9, 1.666789298E9, 1.666789346E9, 1.666789394E9, 1.666789442E9, 1.66678949E9, 1.666789538E9, 1.666789586E9, 1.666789634E9, 1.666789682E9, 1.66678973E9, 1.666789778E9, 1.666789826E9, 1.666789874E9, 1.666789922E9, 1.66678997E9, 1.666790018E9, 1.666790066E9, 1.666790114E9, 1.666790162E9, 1.66679021E9, 1.666790258E9, 1.666790306E9, 1.666790354E9, 1.666790402E9, 1.66679045E9, 1.66679082E9, 1.666791E9, 1.666796677E9, 1.666796725E9, 1.666796773E9, 1.666796821E9, 1.666796869E9, 1.666796917E9, 1.666796965E9, 1.666797013E9, 1.666797061E9, 1.666797109E9, 1.666797157E9, 1.666797205E9, 1.666797253E9, 1.666797301E9, 1.666797349E9, 1.666797397E9, 1.666797445E9, 1.666797493E9, 1.666797541E9, 1.666797589E9, 1.666797637E9, 1.666797685E9, 1.666797733E9, 1.666797781E9, 1.666797829E9, 1.666797877E9, 1.666797925E9, 1.666797973E9, 1.666798021E9, 1.666798069E9, 1.666798117E9, 1.666798165E9, 1.666798213E9, 1.666798261E9, 1.666798309E9, 1.666798357E9, 1.666798405E9, 1.666798453E9, 1.666798501E9, 1.666798549E9, 1.666798597E9, 1.666798645E9, 1.666798693E9, 1.666798741E9, 1.666798789E9, 1.666798837E9, 1.666798885E9, 1.666798933E9, 1.666798981E9, 1.666799029E9, 1.666799077E9, 1.666799125E9, 1.666799173E9, 1.666799221E9, 1.666799269E9, 1.666799317E9, 1.666799365E9, 1.666799413E9, 1.666799461E9, 1.666799509E9, 1.666799557E9, 1.666799605E9, 1.666799653E9, 1.666799701E9, 1.666799749E9, 1.666799797E9, 1.666799845E9, 1.666799893E9, 1.666799941E9, 1.666799989E9, 1.66680036E9, 1.66680054E9, 1.666806348E9, 1.666806396E9, 1.666806444E9, 1.666806492E9, 1.66680654E9, 1.666806588E9, 1.666806636E9, 1.666806684E9, 1.666806732E9, 1.66680678E9, 1.666806828E9, 1.666806876E9, 1.666806924E9, 1.666806972E9, 1.66680702E9, 1.666807068E9, 1.666807116E9, 1.666807164E9, 1.666807212E9, 1.66680726E9, 1.666807308E9, 1.666807356E9, 1.666807404E9, 1.666807452E9, 1.6668075E9, 1.666807548E9, 1.666807596E9, 1.666807644E9, 1.666807692E9, 1.66680774E9, 1.666807788E9, 1.666807836E9, 1.666807884E9, 1.666807932E9, 1.66680798E9, 1.666808028E9, 1.666808076E9, 1.666808124E9, 1.666808172E9, 1.66680822E9, 1.666808268E9, 1.666808316E9, 1.666808364E9, 1.666808412E9, 1.66680846E9, 1.666808508E9, 1.666808556E9, 1.666808604E9, 1.666808652E9, 1.6668087E9, 1.666808748E9, 1.666808796E9, 1.666808844E9, 1.666808892E9, 1.66680894E9, 1.666808988E9, 1.666809036E9, 1.666809084E9, 1.666809132E9, 1.66680918E9, 1.666809228E9, 1.666809276E9, 1.666809324E9, 1.666809372E9, 1.66680942E9, 1.666809468E9, 1.666809516E9, 1.666809564E9, 1.666809612E9, 1.66680966E9, 1.666809708E9, 1.666809756E9, 1.666809804E9, 1.666809852E9, 1.6668099E9, 1.6668102E9, 1.66681038E9, 1.666816285E9, 1.666816333E9, 1.666816381E9, 1.666816429E9, 1.666816477E9, 1.666816525E9, 1.666816573E9, 1.666816621E9, 1.666816669E9, 1.666816717E9, 1.666816765E9, 1.666816813E9, 1.666816861E9, 1.666816909E9, 1.666816957E9, 1.666817005E9, 1.666817053E9, 1.666817101E9, 1.666817149E9, 1.666817197E9, 1.666817245E9, 1.666817293E9, 1.666817341E9, 1.666817389E9, 1.666817437E9, 1.666817485E9, 1.666817533E9, 1.666817581E9, 1.666817629E9, 1.666817677E9, 1.666817725E9, 1.666817773E9, 1.666817821E9, 1.666817869E9, 1.666817917E9, 1.666817965E9, 1.666818013E9, 1.666818061E9, 1.666818109E9, 1.666818157E9, 1.666818205E9, 1.666818253E9, 1.666818301E9, 1.666818349E9, 1.666818397E9, 1.666818445E9, 1.666818493E9, 1.666818541E9, 1.666818589E9, 1.666818637E9, 1.666818685E9, 1.666818733E9, 1.666818781E9, 1.666818829E9, 1.666818877E9, 1.666818925E9, 1.666818973E9, 1.666819021E9, 1.666819069E9, 1.666819117E9, 1.666819165E9, 1.666819213E9, 1.666819261E9, 1.666819309E9, 1.666819357E9, 1.666819405E9, 1.666819453E9, 1.666819501E9, 1.666819549E9, 1.66681992E9, 1.66682004E9, 1.666825842E9, 1.66682589E9, 1.666825938E9, 1.666825986E9, 1.666826034E9, 1.666826082E9, 1.66682613E9, 1.666826178E9, 1.666826226E9, 1.666826274E9, 1.666826322E9, 1.66682637E9, 1.666826418E9, 1.666826466E9, 1.666826514E9, 1.666826562E9, 1.66682661E9, 1.666826658E9, 1.666826706E9, 1.666826754E9, 1.666826802E9, 1.66682685E9, 1.666826898E9, 1.666826946E9, 1.666826994E9, 1.666827042E9, 1.66682709E9, 1.666827138E9, 1.666827186E9, 1.666827234E9, 1.666827282E9, 1.66682733E9, 1.666827378E9, 1.666827426E9, 1.666827474E9, 1.666827522E9, 1.66682757E9, 1.666827618E9, 1.666827666E9, 1.666827714E9, 1.666827762E9, 1.66682781E9, 1.666827858E9, 1.666827906E9, 1.666827954E9, 1.666828002E9, 1.66682805E9, 1.666828098E9, 1.666828146E9, 1.666828194E9, 1.666828242E9, 1.66682829E9, 1.666828338E9, 1.666828386E9, 1.666828434E9, 1.666828482E9, 1.66682853E9, 1.666828578E9, 1.666828626E9, 1.666828674E9, 1.666828722E9, 1.66682877E9, 1.666828818E9, 1.666828866E9, 1.666828914E9, 1.666828962E9, 1.66682901E9, 1.666829058E9, 1.666829106E9, 1.666829154E9, 1.666829202E9, 1.66682925E9, 1.66682958E9, 1.66682976E9, 1.666835651E9, 1.666835699E9, 1.666835747E9, 1.666835795E9, 1.666835843E9, 1.666835891E9, 1.666835939E9, 1.666835987E9, 1.666836035E9, 1.666836083E9, 1.666836131E9, 1.666836179E9, 1.666836227E9, 1.666836275E9, 1.666836323E9, 1.666836371E9, 1.666836419E9, 1.666836467E9, 1.666836515E9, 1.666836563E9, 1.666836611E9, 1.666836659E9, 1.666836707E9, 1.666836755E9, 1.666836803E9, 1.666836851E9, 1.666836899E9, 1.666836947E9, 1.666836995E9, 1.666837043E9, 1.666837091E9, 1.666837139E9, 1.666837187E9, 1.666837235E9, 1.666837283E9, 1.666837331E9, 1.666837379E9, 1.666837427E9, 1.666837475E9, 1.666837523E9, 1.666837571E9, 1.666837619E9, 1.666837667E9, 1.666837715E9, 1.666837763E9, 1.666837811E9, 1.666837859E9, 1.666837907E9, 1.666837955E9, 1.666838003E9, 1.666838051E9, 1.666838099E9, 1.666838147E9, 1.666838195E9, 1.666838243E9, 1.666838291E9, 1.666838339E9, 1.666838387E9, 1.666838435E9, 1.666838483E9, 1.666838531E9, 1.666838579E9, 1.666838627E9, 1.666838675E9, 1.666838723E9, 1.666838771E9, 1.666838819E9, 1.666838867E9, 1.666838915E9, 1.666838963E9, 1.666839011E9, 1.666839059E9, 1.6668393E9, 1.66683948E9, 1.666845277E9, 1.666845325E9, 1.666845373E9, 1.666845421E9, 1.666845469E9, 1.666845517E9, 1.666845565E9, 1.666845613E9, 1.666845661E9, 1.666845709E9, 1.666845757E9, 1.666845805E9, 1.666845853E9, 1.666845901E9, 1.666845949E9, 1.666845997E9, 1.666846045E9, 1.666846093E9, 1.666846141E9, 1.666846189E9, 1.666846237E9, 1.666846285E9, 1.666846333E9, 1.666846381E9, 1.666846429E9, 1.666846477E9, 1.666846525E9, 1.666846573E9, 1.666846621E9, 1.666846669E9, 1.666846717E9, 1.666846765E9, 1.666846813E9, 1.666846861E9, 1.666846909E9, 1.666846957E9, 1.666847005E9, 1.666847053E9, 1.666847101E9, 1.666847149E9, 1.666847197E9, 1.666847245E9, 1.666847293E9, 1.666847341E9, 1.666847389E9, 1.666847437E9, 1.666847485E9, 1.666847533E9, 1.666847581E9, 1.666847629E9, 1.666847677E9, 1.666847725E9, 1.666847773E9, 1.666847821E9, 1.666847869E9, 1.666847917E9, 1.666847965E9, 1.666848013E9, 1.666848061E9, 1.666848109E9, 1.666848157E9, 1.666848205E9, 1.666848253E9, 1.666848301E9, 1.666848349E9, 1.666848397E9, 1.666848445E9, 1.666848493E9, 1.666848541E9, 1.666848589E9, 1.66684896E9, 1.66684914E9, 1.666855042E9, 1.66685509E9, 1.666855138E9, 1.666855186E9, 1.666855234E9, 1.666855282E9, 1.66685533E9, 1.666855378E9, 1.666855426E9, 1.666855474E9, 1.666855522E9, 1.66685557E9, 1.666855618E9, 1.666855666E9, 1.666855714E9, 1.666855762E9, 1.66685581E9, 1.666855858E9, 1.666855906E9, 1.666855954E9, 1.666856002E9, 1.66685605E9, 1.666856098E9, 1.666856146E9, 1.666856194E9, 1.666856242E9, 1.66685629E9, 1.666856338E9, 1.666856386E9, 1.666856434E9, 1.666856482E9, 1.66685653E9, 1.666856578E9, 1.666856626E9, 1.666856674E9, 1.666856722E9, 1.66685677E9, 1.666856818E9, 1.666856866E9, 1.666856914E9, 1.666856962E9, 1.66685701E9, 1.666857058E9, 1.666857106E9, 1.666857154E9, 1.666857202E9, 1.66685725E9, 1.666857298E9, 1.666857346E9, 1.666857394E9, 1.666857442E9, 1.66685749E9, 1.666857538E9, 1.666857586E9, 1.666857634E9, 1.666857682E9, 1.66685773E9, 1.666857778E9, 1.666857826E9, 1.666857874E9, 1.666857922E9, 1.66685797E9, 1.666858018E9, 1.666858066E9, 1.666858114E9, 1.666858162E9, 1.66685821E9, 1.666858258E9, 1.666858306E9, 1.666858354E9, 1.666858402E9, 1.66685845E9, 1.6668588E9, 1.66685898E9, 1.666864666E9, 1.666864714E9, 1.666864762E9, 1.66686481E9, 1.666864858E9, 1.666864906E9, 1.666864954E9, 1.666865002E9, 1.66686505E9, 1.666865098E9, 1.666865146E9, 1.666865194E9, 1.666865242E9, 1.66686529E9, 1.666865338E9, 1.666865386E9, 1.666865434E9, 1.666865482E9, 1.66686553E9, 1.666865578E9, 1.666865626E9, 1.666865674E9, 1.666865722E9, 1.66686577E9, 1.666865818E9, 1.666865866E9, 1.666865914E9, 1.666865962E9, 1.66686601E9, 1.666866058E9, 1.666866106E9, 1.666866154E9, 1.666866202E9, 1.66686625E9, 1.666866298E9, 1.666866346E9, 1.666866394E9, 1.666866442E9, 1.66686649E9, 1.666866538E9, 1.666866586E9, 1.666866634E9, 1.666866682E9, 1.66686673E9, 1.666866778E9, 1.666866826E9, 1.666866874E9, 1.666866922E9, 1.66686697E9, 1.666867018E9, 1.666867066E9, 1.666867114E9, 1.666867162E9, 1.66686721E9, 1.666867258E9, 1.666867306E9, 1.666867354E9, 1.666867402E9, 1.66686745E9, 1.666867498E9, 1.666867546E9, 1.666867594E9, 1.666867642E9, 1.66686769E9, 1.666867738E9, 1.666867786E9, 1.666867834E9, 1.666867882E9, 1.66686793E9, 1.66686828E9, 1.66686846E9, 1.666874535E9, 1.666874583E9, 1.666874631E9, 1.666874679E9, 1.666874727E9, 1.666874775E9, 1.666874823E9, 1.666874871E9, 1.666874919E9, 1.666874967E9, 1.666875015E9, 1.666875063E9, 1.666875111E9, 1.666875159E9, 1.666875207E9, 1.666875255E9, 1.666875303E9, 1.666875351E9, 1.666875399E9, 1.666875447E9, 1.666875495E9, 1.666875543E9, 1.666875591E9, 1.666875639E9, 1.666875687E9, 1.666875735E9, 1.666875783E9, 1.666875831E9, 1.666875879E9, 1.666875927E9, 1.666875975E9, 1.666876023E9, 1.666876071E9, 1.666876119E9, 1.666876167E9, 1.666876215E9, 1.666876263E9, 1.666876311E9, 1.666876359E9, 1.666876407E9, 1.666876455E9, 1.666876503E9, 1.666876551E9, 1.666876599E9, 1.666876647E9, 1.666876695E9, 1.666876743E9, 1.666876791E9, 1.666876839E9, 1.666876887E9, 1.666876935E9, 1.666876983E9, 1.666877031E9, 1.666877079E9, 1.666877127E9, 1.666877175E9, 1.666877223E9, 1.666877271E9, 1.666877319E9, 1.666877367E9, 1.666877415E9, 1.666877463E9, 1.666877511E9, 1.666877559E9, 1.666877607E9, 1.666877655E9, 1.666877703E9, 1.666877751E9, 1.666877799E9, 1.666877847E9, 1.666877895E9, 1.666877943E9, 1.666877991E9, 1.666878039E9, 1.66687842E9, 1.6668786E9, 1.666884676E9, 1.666884724E9, 1.666884772E9, 1.66688482E9, 1.666884868E9, 1.666884916E9, 1.666884964E9, 1.666885012E9, 1.66688506E9, 1.666885108E9, 1.666885156E9, 1.666885204E9, 1.666885252E9, 1.6668853E9, 1.666885348E9, 1.666885396E9, 1.666885444E9, 1.666885492E9, 1.66688554E9, 1.666885588E9, 1.666885636E9, 1.666885684E9, 1.666885732E9, 1.66688578E9, 1.666885828E9, 1.666885876E9, 1.666885924E9, 1.666885972E9, 1.66688602E9, 1.666886068E9, 1.666886116E9, 1.666886164E9, 1.666886212E9, 1.66688626E9, 1.666886308E9, 1.666886356E9, 1.666886404E9, 1.666886452E9, 1.6668865E9, 1.666886548E9, 1.666886596E9, 1.666886644E9, 1.666886692E9, 1.66688674E9, 1.666886788E9, 1.666886836E9, 1.666886884E9, 1.666886932E9, 1.66688698E9, 1.666887028E9, 1.666887076E9, 1.666887124E9, 1.666887172E9, 1.66688722E9, 1.666887268E9, 1.666887316E9, 1.666887364E9, 1.666887412E9, 1.66688746E9, 1.666887508E9, 1.666887556E9, 1.666887604E9, 1.666887652E9, 1.6668877E9, 1.666887748E9, 1.666887796E9, 1.666887844E9, 1.666887892E9, 1.66688794E9, 1.66688832E9, 1.6668885E9, 1.666894379E9, 1.666894427E9, 1.666894475E9, 1.666894523E9, 1.666894571E9, 1.666894619E9, 1.666894667E9, 1.666894715E9, 1.666894763E9, 1.666894811E9, 1.666894859E9, 1.666894907E9, 1.666894955E9, 1.666895003E9, 1.666895051E9, 1.666895099E9, 1.666895147E9, 1.666895195E9, 1.666895243E9, 1.666895291E9, 1.666895339E9, 1.666895387E9, 1.666895435E9, 1.666895483E9, 1.666895531E9, 1.666895579E9, 1.666895627E9, 1.666895675E9, 1.666895723E9, 1.666895771E9, 1.666895819E9, 1.666895867E9, 1.666895915E9, 1.666895963E9, 1.666896011E9, 1.666896059E9, 1.666896107E9, 1.666896155E9, 1.666896203E9, 1.666896251E9, 1.666896299E9, 1.666896347E9, 1.666896395E9, 1.666896443E9, 1.666896491E9, 1.666896539E9, 1.666896587E9, 1.666896635E9, 1.666896683E9, 1.666896731E9, 1.666896779E9, 1.666896827E9, 1.666896875E9, 1.666896923E9, 1.666896971E9, 1.666897019E9, 1.666897067E9, 1.666897115E9, 1.666897163E9, 1.666897211E9, 1.666897259E9, 1.666897307E9, 1.666897355E9, 1.666897403E9, 1.666897451E9, 1.666897499E9, 1.666897547E9, 1.666897595E9, 1.666897643E9, 1.666897691E9, 1.666897739E9, 1.66689804E9, 1.66689822E9, 1.666903864E9, 1.666903912E9, 1.66690396E9, 1.666904008E9, 1.666904056E9, 1.666904104E9, 1.666904152E9, 1.6669042E9, 1.666904248E9, 1.666904296E9, 1.666904344E9, 1.666904392E9, 1.66690444E9, 1.666904488E9, 1.666904536E9, 1.666904584E9, 1.666904632E9, 1.66690468E9, 1.666904728E9, 1.666904776E9, 1.666904824E9, 1.666904872E9, 1.66690492E9, 1.666904968E9, 1.666905016E9, 1.666905064E9, 1.666905112E9, 1.66690516E9, 1.666905208E9, 1.666905256E9, 1.666905304E9, 1.666905352E9, 1.6669054E9, 1.666905448E9, 1.666905496E9, 1.666905544E9, 1.666905592E9, 1.66690564E9, 1.666905688E9, 1.666905736E9, 1.666905784E9, 1.666905832E9, 1.66690588E9, 1.666905928E9, 1.666905976E9, 1.666906024E9, 1.666906072E9, 1.66690612E9, 1.666906168E9, 1.666906216E9, 1.666906264E9, 1.666906312E9, 1.66690636E9, 1.666906408E9, 1.666906456E9, 1.666906504E9, 1.666906552E9, 1.6669066E9, 1.666906648E9, 1.666906696E9, 1.666906744E9, 1.666906792E9, 1.66690684E9, 1.666906888E9, 1.666906936E9, 1.666906984E9, 1.666907032E9, 1.66690708E9, 1.6669074E9, 1.66690758E9, 1.666913495E9, 1.666913543E9, 1.666913591E9, 1.666913639E9, 1.666913687E9, 1.666913735E9, 1.666913783E9, 1.666913831E9, 1.666913879E9, 1.666913927E9, 1.666913975E9, 1.666914023E9, 1.666914071E9, 1.666914119E9, 1.666914167E9, 1.666914215E9, 1.666914263E9, 1.666914311E9, 1.666914359E9, 1.666914407E9, 1.666914455E9, 1.666914503E9, 1.666914551E9, 1.666914599E9, 1.666914647E9, 1.666914695E9, 1.666914743E9, 1.666914791E9, 1.666914839E9, 1.666914887E9, 1.666914935E9, 1.666914983E9, 1.666915031E9, 1.666915079E9, 1.666915127E9, 1.666915175E9, 1.666915223E9, 1.666915271E9, 1.666915319E9, 1.666915367E9, 1.666915415E9, 1.666915463E9, 1.666915511E9, 1.666915559E9, 1.666915607E9, 1.666915655E9, 1.666915703E9, 1.666915751E9, 1.666915799E9, 1.666915847E9, 1.666915895E9, 1.666915943E9, 1.666915991E9, 1.666916039E9, 1.666916087E9, 1.666916135E9, 1.666916183E9, 1.666916231E9, 1.666916279E9, 1.666916327E9, 1.666916375E9, 1.666916423E9, 1.666916471E9, 1.666916519E9, 1.666916567E9, 1.666916615E9, 1.666916663E9, 1.666916711E9, 1.666916759E9, 1.66691712E9, 1.6669173E9, 1.66692313E9, 1.666923178E9, 1.666923226E9, 1.666923274E9, 1.666923322E9, 1.66692337E9, 1.666923418E9, 1.666923466E9, 1.666923514E9, 1.666923562E9, 1.66692361E9, 1.666923658E9, 1.666923706E9, 1.666923754E9, 1.666923802E9, 1.66692385E9, 1.666923898E9, 1.666923946E9, 1.666923994E9, 1.666924042E9, 1.66692409E9, 1.666924138E9, 1.666924186E9, 1.666924234E9, 1.666924282E9, 1.66692433E9, 1.666924378E9, 1.666924426E9, 1.666924474E9, 1.666924522E9, 1.66692457E9, 1.666924618E9, 1.666924666E9, 1.666924714E9, 1.666924762E9, 1.66692481E9, 1.666924858E9, 1.666924906E9, 1.666924954E9, 1.666925002E9, 1.66692505E9, 1.666925098E9, 1.666925146E9, 1.666925194E9, 1.666925242E9, 1.66692529E9, 1.666925338E9, 1.666925386E9, 1.666925434E9, 1.666925482E9, 1.66692553E9, 1.666925578E9, 1.666925626E9, 1.666925674E9, 1.666925722E9, 1.66692577E9, 1.666925818E9, 1.666925866E9, 1.666925914E9, 1.666925962E9, 1.66692601E9, 1.666926058E9, 1.666926106E9, 1.666926154E9, 1.666926202E9, 1.66692625E9, 1.666926298E9, 1.666926346E9, 1.666926394E9, 1.666926442E9, 1.66692649E9, 1.66692678E9, 1.66692696E9, 1.666932963E9, 1.666933011E9, 1.666933059E9, 1.666933107E9, 1.666933155E9, 1.666933203E9, 1.666933251E9, 1.666933299E9, 1.666933347E9, 1.666933395E9, 1.666933443E9, 1.666933491E9, 1.666933539E9, 1.666933587E9, 1.666933635E9, 1.666933683E9, 1.666933731E9, 1.666933779E9, 1.666933827E9, 1.666933875E9, 1.666933923E9, 1.666933971E9, 1.666934019E9, 1.666934067E9, 1.666934115E9, 1.666934163E9, 1.666934211E9, 1.666934259E9, 1.666934307E9, 1.666934355E9, 1.666934403E9, 1.666934451E9, 1.666934499E9, 1.666934547E9, 1.666934595E9, 1.666934643E9, 1.666934691E9, 1.666934739E9, 1.666934787E9, 1.666934835E9, 1.666934883E9, 1.666934931E9, 1.666934979E9, 1.666935027E9, 1.666935075E9, 1.666935123E9, 1.666935171E9, 1.666935219E9, 1.666935267E9, 1.666935315E9, 1.666935363E9, 1.666935411E9, 1.666935459E9, 1.666935507E9, 1.666935555E9, 1.666935603E9, 1.666935651E9, 1.666935699E9, 1.666935747E9, 1.666935795E9, 1.666935843E9, 1.666935891E9, 1.666935939E9, 1.666935987E9, 1.666936035E9, 1.666936083E9, 1.666936131E9, 1.666936179E9, 1.666936227E9, 1.666936275E9, 1.666936323E9, 1.666936371E9, 1.666936419E9, 1.666936467E9, 1.666936515E9, 1.666936563E9, 1.666936611E9, 1.666936659E9, 1.66693704E9, 1.66693722E9, 1.666943072E9, 1.66694312E9, 1.666943168E9, 1.666943216E9, 1.666943264E9, 1.666943312E9, 1.66694336E9, 1.666943408E9, 1.666943456E9, 1.666943504E9, 1.666943552E9, 1.6669436E9, 1.666943648E9, 1.666943696E9, 1.666943744E9, 1.666943792E9, 1.66694384E9, 1.666943888E9, 1.666943936E9, 1.666943984E9, 1.666944032E9, 1.66694408E9, 1.666944128E9, 1.666944176E9, 1.666944224E9, 1.666944272E9, 1.66694432E9, 1.666944368E9, 1.666944416E9, 1.666944464E9, 1.666944512E9, 1.66694456E9, 1.666944608E9, 1.666944656E9, 1.666944704E9, 1.666944752E9, 1.6669448E9, 1.666944848E9, 1.666944896E9, 1.666944944E9, 1.666944992E9, 1.66694504E9, 1.666945088E9, 1.666945136E9, 1.666945184E9, 1.666945232E9, 1.66694528E9, 1.666945328E9, 1.666945376E9, 1.666945424E9, 1.666945472E9, 1.66694552E9, 1.666945568E9, 1.666945616E9, 1.666945664E9, 1.666945712E9, 1.66694576E9, 1.666945808E9, 1.666945856E9, 1.666945904E9, 1.666945952E9, 1.666946E9, 1.666946048E9, 1.666946096E9, 1.666946144E9, 1.666946192E9, 1.66694624E9, 1.66694652E9, 1.6669467E9, 1.666952479E9, 1.666952527E9, 1.666952575E9, 1.666952623E9, 1.666952671E9, 1.666952719E9, 1.666952767E9, 1.666952815E9, 1.666952863E9, 1.666952911E9, 1.666952959E9, 1.666953007E9, 1.666953055E9, 1.666953103E9, 1.666953151E9, 1.666953199E9, 1.666953247E9, 1.666953295E9, 1.666953343E9, 1.666953391E9, 1.666953439E9, 1.666953487E9, 1.666953535E9, 1.666953583E9, 1.666953631E9, 1.666953679E9, 1.666953727E9, 1.666953775E9, 1.666953823E9, 1.666953871E9, 1.666953919E9, 1.666953967E9, 1.666954015E9, 1.666954063E9, 1.666954111E9, 1.666954159E9, 1.666954207E9, 1.666954255E9, 1.666954303E9, 1.666954351E9, 1.666954399E9, 1.666954447E9, 1.666954495E9, 1.666954543E9, 1.666954591E9, 1.666954639E9, 1.666954687E9, 1.666954735E9, 1.666954783E9, 1.666954831E9, 1.666954879E9, 1.666954927E9, 1.666954975E9, 1.666955023E9, 1.666955071E9, 1.666955119E9, 1.666955167E9, 1.666955215E9, 1.666955263E9, 1.666955311E9, 1.666955359E9, 1.666955407E9, 1.666955455E9, 1.666955503E9, 1.666955551E9, 1.666955599E9, 1.666955647E9, 1.666955695E9, 1.666955743E9, 1.666955791E9, 1.666955839E9, 1.66695612E9, 1.66695636E9, 1.666962244E9, 1.666962292E9, 1.66696234E9, 1.666962388E9, 1.666962436E9, 1.666962484E9, 1.666962532E9, 1.66696258E9, 1.666962628E9, 1.666962676E9, 1.666962724E9, 1.666962772E9, 1.66696282E9, 1.666962868E9, 1.666962916E9, 1.666962964E9, 1.666963012E9, 1.66696306E9, 1.666963108E9, 1.666963156E9, 1.666963204E9, 1.666963252E9, 1.6669633E9, 1.666963348E9, 1.666963396E9, 1.666963444E9, 1.666963492E9, 1.66696354E9, 1.666963588E9, 1.666963636E9, 1.666963684E9, 1.666963732E9, 1.66696378E9, 1.666963828E9, 1.666963876E9, 1.666963924E9, 1.666963972E9, 1.66696402E9, 1.666964068E9, 1.666964116E9, 1.666964164E9, 1.666964212E9, 1.66696426E9, 1.666964308E9, 1.666964356E9, 1.666964404E9, 1.666964452E9, 1.6669645E9, 1.666964548E9, 1.666964596E9, 1.666964644E9, 1.666964692E9, 1.66696474E9, 1.666964788E9, 1.666964836E9, 1.666964884E9, 1.666964932E9, 1.66696498E9, 1.666965028E9, 1.666965076E9, 1.666965124E9, 1.666965172E9, 1.66696522E9, 1.666965268E9, 1.666965316E9, 1.666965364E9, 1.666965412E9, 1.66696546E9, 1.66696578E9, 1.66696596E9, 1.66697179E9, 1.666971838E9, 1.666971886E9, 1.666971934E9, 1.666971982E9, 1.66697203E9, 1.666972078E9, 1.666972126E9, 1.666972174E9, 1.666972222E9, 1.66697227E9, 1.666972318E9, 1.666972366E9, 1.666972414E9, 1.666972462E9, 1.66697251E9, 1.666972558E9, 1.666972606E9, 1.666972654E9, 1.666972702E9, 1.66697275E9, 1.666972798E9, 1.666972846E9, 1.666972894E9, 1.666972942E9, 1.66697299E9, 1.666973038E9, 1.666973086E9, 1.666973134E9, 1.666973182E9, 1.66697323E9, 1.666973278E9, 1.666973326E9, 1.666973374E9, 1.666973422E9, 1.66697347E9, 1.666973518E9, 1.666973566E9, 1.666973614E9, 1.666973662E9, 1.66697371E9, 1.666973758E9, 1.666973806E9, 1.666973854E9, 1.666973902E9, 1.66697395E9, 1.666973998E9, 1.666974046E9, 1.666974094E9, 1.666974142E9, 1.66697419E9, 1.666974238E9, 1.666974286E9, 1.666974334E9, 1.666974382E9, 1.66697443E9, 1.666974478E9, 1.666974526E9, 1.666974574E9, 1.666974622E9, 1.66697467E9, 1.666974718E9, 1.666974766E9, 1.666974814E9, 1.666974862E9, 1.66697491E9, 1.666974958E9, 1.666975006E9, 1.666975054E9, 1.666975102E9, 1.66697515E9, 1.66697544E9, 1.66697562E9, 1.66698141E9, 1.666981458E9, 1.666981506E9, 1.666981554E9, 1.666981602E9, 1.66698165E9, 1.666981698E9, 1.666981746E9, 1.666981794E9, 1.666981842E9, 1.66698189E9, 1.666981938E9, 1.666981986E9, 1.666982034E9, 1.666982082E9, 1.66698213E9, 1.666982178E9, 1.666982226E9, 1.666982274E9, 1.666982322E9, 1.66698237E9, 1.666982418E9, 1.666982466E9, 1.666982514E9, 1.666982562E9, 1.66698261E9, 1.666982658E9, 1.666982706E9, 1.666982754E9, 1.666982802E9, 1.66698285E9, 1.666982898E9, 1.666982946E9, 1.666982994E9, 1.666983042E9, 1.66698309E9, 1.666983138E9, 1.666983186E9, 1.666983234E9, 1.666983282E9, 1.66698333E9, 1.666983378E9, 1.666983426E9, 1.666983474E9, 1.666983522E9, 1.66698357E9, 1.666983618E9, 1.666983666E9, 1.666983714E9, 1.666983762E9, 1.66698381E9, 1.666983858E9, 1.666983906E9, 1.666983954E9, 1.666984002E9, 1.66698405E9, 1.666984098E9, 1.666984146E9, 1.666984194E9, 1.666984242E9, 1.66698429E9, 1.666984338E9, 1.666984386E9, 1.666984434E9, 1.666984482E9, 1.66698453E9, 1.666984578E9, 1.666984626E9, 1.666984674E9, 1.666984722E9, 1.66698477E9, 1.666984818E9, 1.666984866E9, 1.666984914E9, 1.666984962E9, 1.66698501E9, 1.66698534E9, 1.66698552E9, 1.666991353E9, 1.666991401E9, 1.666991449E9, 1.666991497E9, 1.666991545E9, 1.666991593E9, 1.666991641E9, 1.666991689E9, 1.666991737E9, 1.666991785E9, 1.666991833E9, 1.666991881E9, 1.666991929E9, 1.666991977E9, 1.666992025E9, 1.666992073E9, 1.666992121E9, 1.666992169E9, 1.666992217E9, 1.666992265E9, 1.666992313E9, 1.666992361E9, 1.666992409E9, 1.666992457E9, 1.666992505E9, 1.666992553E9, 1.666992601E9, 1.666992649E9, 1.666992697E9, 1.666992745E9, 1.666992793E9, 1.666992841E9, 1.666992889E9, 1.666992937E9, 1.666992985E9, 1.666993033E9, 1.666993081E9, 1.666993129E9, 1.666993177E9, 1.666993225E9, 1.666993273E9, 1.666993321E9, 1.666993369E9, 1.666993417E9, 1.666993465E9, 1.666993513E9, 1.666993561E9, 1.666993609E9, 1.666993657E9, 1.666993705E9, 1.666993753E9, 1.666993801E9, 1.666993849E9, 1.666993897E9, 1.666993945E9, 1.666993993E9, 1.666994041E9, 1.666994089E9, 1.666994137E9, 1.666994185E9, 1.666994233E9, 1.666994281E9, 1.666994329E9, 1.666994377E9, 1.666994425E9, 1.666994473E9, 1.666994521E9, 1.666994569E9, 1.66699488E9, 1.66699506E9, 1.667000929E9, 1.667000977E9, 1.667001025E9, 1.667001073E9, 1.667001121E9, 1.667001169E9, 1.667001217E9, 1.667001265E9, 1.667001313E9, 1.667001361E9, 1.667001409E9, 1.667001457E9, 1.667001505E9, 1.667001553E9, 1.667001601E9, 1.667001649E9, 1.667001697E9, 1.667001745E9, 1.667001793E9, 1.667001841E9, 1.667001889E9, 1.667001937E9, 1.667001985E9, 1.667002033E9, 1.667002081E9, 1.667002129E9, 1.667002177E9, 1.667002225E9, 1.667002273E9, 1.667002321E9, 1.667002369E9, 1.667002417E9, 1.667002465E9, 1.667002513E9, 1.667002561E9, 1.667002609E9, 1.667002657E9, 1.667002705E9, 1.667002753E9, 1.667002801E9, 1.667002849E9, 1.667002897E9, 1.667002945E9, 1.667002993E9, 1.667003041E9, 1.667003089E9, 1.667003137E9, 1.667003185E9, 1.667003233E9, 1.667003281E9, 1.667003329E9, 1.667003377E9, 1.667003425E9, 1.667003473E9, 1.667003521E9, 1.667003569E9, 1.667003617E9, 1.667003665E9, 1.667003713E9, 1.667003761E9, 1.667003809E9, 1.667003857E9, 1.667003905E9, 1.667003953E9, 1.667004001E9, 1.667004049E9, 1.66700436E9, 1.66700454E9, 1.66701037E9, 1.667010418E9, 1.667010466E9, 1.667010514E9, 1.667010562E9, 1.66701061E9, 1.667010658E9, 1.667010706E9, 1.667010754E9, 1.667010802E9, 1.66701085E9, 1.667010898E9, 1.667010946E9, 1.667010994E9, 1.667011042E9, 1.66701109E9, 1.667011138E9, 1.667011186E9, 1.667011234E9, 1.667011282E9, 1.66701133E9, 1.667011378E9, 1.667011426E9, 1.667011474E9, 1.667011522E9, 1.66701157E9, 1.667011618E9, 1.667011666E9, 1.667011714E9, 1.667011762E9, 1.66701181E9, 1.667011858E9, 1.667011906E9, 1.667011954E9, 1.667012002E9, 1.66701205E9, 1.667012098E9, 1.667012146E9, 1.667012194E9, 1.667012242E9, 1.66701229E9, 1.667012338E9, 1.667012386E9, 1.667012434E9, 1.667012482E9, 1.66701253E9, 1.667012578E9, 1.667012626E9, 1.667012674E9, 1.667012722E9, 1.66701277E9, 1.667012818E9, 1.667012866E9, 1.667012914E9, 1.667012962E9, 1.66701301E9, 1.667013058E9, 1.667013106E9, 1.667013154E9, 1.667013202E9, 1.66701325E9, 1.667013298E9, 1.667013346E9, 1.667013394E9, 1.667013442E9, 1.66701349E9, 1.667013538E9, 1.667013586E9, 1.667013634E9, 1.667013682E9, 1.66701373E9, 1.66701402E9, 1.6670142E9, 1.667020061E9, 1.667020109E9, 1.667020157E9, 1.667020205E9, 1.667020253E9, 1.667020301E9, 1.667020349E9, 1.667020397E9, 1.667020445E9, 1.667020493E9, 1.667020541E9, 1.667020589E9, 1.667020637E9, 1.667020685E9, 1.667020733E9, 1.667020781E9, 1.667020829E9, 1.667020877E9, 1.667020925E9, 1.667020973E9, 1.667021021E9, 1.667021069E9, 1.667021117E9, 1.667021165E9, 1.667021213E9, 1.667021261E9, 1.667021309E9, 1.667021357E9, 1.667021405E9, 1.667021453E9, 1.667021501E9, 1.667021549E9, 1.667021597E9, 1.667021645E9, 1.667021693E9, 1.667021741E9, 1.667021789E9, 1.667021837E9, 1.667021885E9, 1.667021933E9, 1.667021981E9, 1.667022029E9, 1.667022077E9, 1.667022125E9, 1.667022173E9, 1.667022221E9, 1.667022269E9, 1.667022317E9, 1.667022365E9, 1.667022413E9, 1.667022461E9, 1.667022509E9, 1.667022557E9, 1.667022605E9, 1.667022653E9, 1.667022701E9, 1.667022749E9, 1.667022797E9, 1.667022845E9, 1.667022893E9, 1.667022941E9, 1.667022989E9, 1.667023037E9, 1.667023085E9, 1.667023133E9, 1.667023181E9, 1.667023229E9, 1.667023277E9, 1.667023325E9, 1.667023373E9, 1.667023421E9, 1.667023469E9, 1.66702374E9, 1.66702392E9, 1.667029858E9, 1.667029906E9, 1.667029954E9, 1.667030002E9, 1.66703005E9, 1.667030098E9, 1.667030146E9, 1.667030194E9, 1.667030242E9, 1.66703029E9, 1.667030338E9, 1.667030386E9, 1.667030434E9, 1.667030482E9, 1.66703053E9, 1.667030578E9, 1.667030626E9, 1.667030674E9, 1.667030722E9, 1.66703077E9, 1.667030818E9, 1.667030866E9, 1.667030914E9, 1.667030962E9, 1.66703101E9, 1.667031058E9, 1.667031106E9, 1.667031154E9, 1.667031202E9, 1.66703125E9, 1.667031298E9, 1.667031346E9, 1.667031394E9, 1.667031442E9, 1.66703149E9, 1.667031538E9, 1.667031586E9, 1.667031634E9, 1.667031682E9, 1.66703173E9, 1.667031778E9, 1.667031826E9, 1.667031874E9, 1.667031922E9, 1.66703197E9, 1.667032018E9, 1.667032066E9, 1.667032114E9, 1.667032162E9, 1.66703221E9, 1.667032258E9, 1.667032306E9, 1.667032354E9, 1.667032402E9, 1.66703245E9, 1.667032498E9, 1.667032546E9, 1.667032594E9, 1.667032642E9, 1.66703269E9, 1.667032738E9, 1.667032786E9, 1.667032834E9, 1.667032882E9, 1.66703293E9, 1.667032978E9, 1.667033026E9, 1.667033074E9, 1.667033122E9, 1.66703317E9, 1.66703346E9, 1.66703364E9, 1.667039345E9, 1.667039393E9, 1.667039441E9, 1.667039489E9, 1.667039537E9, 1.667039585E9, 1.667039633E9, 1.667039681E9, 1.667039729E9, 1.667039777E9, 1.667039825E9, 1.667039873E9, 1.667039921E9, 1.667039969E9, 1.667040017E9, 1.667040065E9, 1.667040113E9, 1.667040161E9, 1.667040209E9, 1.667040257E9, 1.667040305E9, 1.667040353E9, 1.667040401E9, 1.667040449E9, 1.667040497E9, 1.667040545E9, 1.667040593E9, 1.667040641E9, 1.667040689E9, 1.667040737E9, 1.667040785E9, 1.667040833E9, 1.667040881E9, 1.667040929E9, 1.667040977E9, 1.667041025E9, 1.667041073E9, 1.667041121E9, 1.667041169E9, 1.667041217E9, 1.667041265E9, 1.667041313E9, 1.667041361E9, 1.667041409E9, 1.667041457E9, 1.667041505E9, 1.667041553E9, 1.667041601E9, 1.667041649E9, 1.667041697E9, 1.667041745E9, 1.667041793E9, 1.667041841E9, 1.667041889E9, 1.667041937E9, 1.667041985E9, 1.667042033E9, 1.667042081E9, 1.667042129E9, 1.667042177E9, 1.667042225E9, 1.667042273E9, 1.667042321E9, 1.667042369E9, 1.667042417E9, 1.667042465E9, 1.667042513E9, 1.667042561E9, 1.667042609E9, 1.667042657E9, 1.667042705E9, 1.667042753E9, 1.667042801E9, 1.667042849E9, 1.66704312E9, 1.6670433E9, 1.667049349E9, 1.667049397E9, 1.667049445E9, 1.667049493E9, 1.667049541E9, 1.667049589E9, 1.667049637E9, 1.667049685E9, 1.667049733E9, 1.667049781E9, 1.667049829E9, 1.667049877E9, 1.667049925E9, 1.667049973E9, 1.667050021E9, 1.667050069E9, 1.667050117E9, 1.667050165E9, 1.667050213E9, 1.667050261E9, 1.667050309E9, 1.667050357E9, 1.667050405E9, 1.667050453E9, 1.667050501E9, 1.667050549E9, 1.667050597E9, 1.667050645E9, 1.667050693E9, 1.667050741E9, 1.667050789E9, 1.667050837E9, 1.667050885E9, 1.667050933E9, 1.667050981E9, 1.667051029E9, 1.667051077E9, 1.667051125E9, 1.667051173E9, 1.667051221E9, 1.667051269E9, 1.667051317E9, 1.667051365E9, 1.667051413E9, 1.667051461E9, 1.667051509E9, 1.667051557E9, 1.667051605E9, 1.667051653E9, 1.667051701E9, 1.667051749E9, 1.667051797E9, 1.667051845E9, 1.667051893E9, 1.667051941E9, 1.667051989E9, 1.667052037E9, 1.667052085E9, 1.667052133E9, 1.667052181E9, 1.667052229E9, 1.667052277E9, 1.667052325E9, 1.667052373E9, 1.667052421E9, 1.667052469E9, 1.66705278E9, 1.66705296E9, 1.667058677E9, 1.667058725E9, 1.667058773E9, 1.667058821E9, 1.667058869E9, 1.667058917E9, 1.667058965E9, 1.667059013E9, 1.667059061E9, 1.667059109E9, 1.667059157E9, 1.667059205E9, 1.667059253E9, 1.667059301E9, 1.667059349E9, 1.667059397E9, 1.667059445E9, 1.667059493E9, 1.667059541E9, 1.667059589E9, 1.667059637E9, 1.667059685E9, 1.667059733E9, 1.667059781E9, 1.667059829E9, 1.667059877E9, 1.667059925E9, 1.667059973E9, 1.667060021E9, 1.667060069E9, 1.667060117E9, 1.667060165E9, 1.667060213E9, 1.667060261E9, 1.667060309E9, 1.667060357E9, 1.667060405E9, 1.667060453E9, 1.667060501E9, 1.667060549E9, 1.667060597E9, 1.667060645E9, 1.667060693E9, 1.667060741E9, 1.667060789E9, 1.667060837E9, 1.667060885E9, 1.667060933E9, 1.667060981E9, 1.667061029E9, 1.667061077E9, 1.667061125E9, 1.667061173E9, 1.667061221E9, 1.667061269E9, 1.667061317E9, 1.667061365E9, 1.667061413E9, 1.667061461E9, 1.667061509E9, 1.667061557E9, 1.667061605E9, 1.667061653E9, 1.667061701E9, 1.667061749E9, 1.667061797E9, 1.667061845E9, 1.667061893E9, 1.667061941E9, 1.667061989E9, 1.66706226E9, 1.66706244E9, 1.667068477E9, 1.667068525E9, 1.667068573E9, 1.667068621E9, 1.667068669E9, 1.667068717E9, 1.667068765E9, 1.667068813E9, 1.667068861E9, 1.667068909E9, 1.667068957E9, 1.667069005E9, 1.667069053E9, 1.667069101E9, 1.667069149E9, 1.667069197E9, 1.667069245E9, 1.667069293E9, 1.667069341E9, 1.667069389E9, 1.667069437E9, 1.667069485E9, 1.667069533E9, 1.667069581E9, 1.667069629E9, 1.667069677E9, 1.667069725E9, 1.667069773E9, 1.667069821E9, 1.667069869E9, 1.667069917E9, 1.667069965E9, 1.667070013E9, 1.667070061E9, 1.667070109E9, 1.667070157E9, 1.667070205E9, 1.667070253E9, 1.667070301E9, 1.667070349E9, 1.667070397E9, 1.667070445E9, 1.667070493E9, 1.667070541E9, 1.667070589E9, 1.667070637E9, 1.667070685E9, 1.667070733E9, 1.667070781E9, 1.667070829E9, 1.667070877E9, 1.667070925E9, 1.667070973E9, 1.667071021E9, 1.667071069E9, 1.667071117E9, 1.667071165E9, 1.667071213E9, 1.667071261E9, 1.667071309E9, 1.667071357E9, 1.667071405E9, 1.667071453E9, 1.667071501E9, 1.667071549E9, 1.667071597E9, 1.667071645E9, 1.667071693E9, 1.667071741E9, 1.667071789E9, 1.667071837E9, 1.667071885E9, 1.667071933E9, 1.667071981E9, 1.667072029E9, 1.667072077E9, 1.667072125E9, 1.667072173E9, 1.667072221E9, 1.667072269E9, 1.66707252E9, 1.6670727E9, 1.667078392E9, 1.66707844E9, 1.667078488E9, 1.667078536E9, 1.667078584E9, 1.667078632E9, 1.66707868E9, 1.667078728E9, 1.667078776E9, 1.667078824E9, 1.667078872E9, 1.66707892E9, 1.667078968E9, 1.667079016E9, 1.667079064E9, 1.667079112E9, 1.66707916E9, 1.667079208E9, 1.667079256E9, 1.667079304E9, 1.667079352E9, 1.6670794E9, 1.667079448E9, 1.667079496E9, 1.667079544E9, 1.667079592E9, 1.66707964E9, 1.667079688E9, 1.667079736E9, 1.667079784E9, 1.667079832E9, 1.66707988E9, 1.667079928E9, 1.667079976E9, 1.667080024E9, 1.667080072E9, 1.66708012E9, 1.667080168E9, 1.667080216E9, 1.667080264E9, 1.667080312E9, 1.66708036E9, 1.667080408E9, 1.667080456E9, 1.667080504E9, 1.667080552E9, 1.6670806E9, 1.667080648E9, 1.667080696E9, 1.667080744E9, 1.667080792E9, 1.66708084E9, 1.667080888E9, 1.667080936E9, 1.667080984E9, 1.667081032E9, 1.66708108E9, 1.667081128E9, 1.667081176E9, 1.667081224E9, 1.667081272E9, 1.66708132E9, 1.667081368E9, 1.667081416E9, 1.667081464E9, 1.667081512E9, 1.66708156E9, 1.66708188E9, 1.66708206E9, 1.66708787E9, 1.667087918E9, 1.667087966E9, 1.667088014E9, 1.667088062E9, 1.66708811E9, 1.667088158E9, 1.667088206E9, 1.667088254E9, 1.667088302E9, 1.66708835E9, 1.667088398E9, 1.667088446E9, 1.667088494E9, 1.667088542E9, 1.66708859E9, 1.667088638E9, 1.667088686E9, 1.667088734E9, 1.667088782E9, 1.66708883E9, 1.667088878E9, 1.667088926E9, 1.667088974E9, 1.667089022E9, 1.66708907E9, 1.667089118E9, 1.667089166E9, 1.667089214E9, 1.667089262E9, 1.66708931E9, 1.667089358E9, 1.667089406E9, 1.667089454E9, 1.667089502E9, 1.66708955E9, 1.667089598E9, 1.667089646E9, 1.667089694E9, 1.667089742E9, 1.66708979E9, 1.667089838E9, 1.667089886E9, 1.667089934E9, 1.667089982E9, 1.66709003E9, 1.667090078E9, 1.667090126E9, 1.667090174E9, 1.667090222E9, 1.66709027E9, 1.667090318E9, 1.667090366E9, 1.667090414E9, 1.667090462E9, 1.66709051E9, 1.667090558E9, 1.667090606E9, 1.667090654E9, 1.667090702E9, 1.66709075E9, 1.667090798E9, 1.667090846E9, 1.667090894E9, 1.667090942E9, 1.66709099E9, 1.667091038E9, 1.667091086E9, 1.667091134E9, 1.667091182E9, 1.66709123E9, 1.66709154E9, 1.66709172E9, 1.667097482E9, 1.66709753E9, 1.667097578E9, 1.667097626E9, 1.667097674E9, 1.667097722E9, 1.66709777E9, 1.667097818E9, 1.667097866E9, 1.667097914E9, 1.667097962E9, 1.66709801E9, 1.667098058E9, 1.667098106E9, 1.667098154E9, 1.667098202E9, 1.66709825E9, 1.667098298E9, 1.667098346E9, 1.667098394E9, 1.667098442E9, 1.66709849E9, 1.667098538E9, 1.667098586E9, 1.667098634E9, 1.667098682E9, 1.66709873E9, 1.667098778E9, 1.667098826E9, 1.667098874E9, 1.667098922E9, 1.66709897E9, 1.667099018E9, 1.667099066E9, 1.667099114E9, 1.667099162E9, 1.66709921E9, 1.667099258E9, 1.667099306E9, 1.667099354E9, 1.667099402E9, 1.66709945E9, 1.667099498E9, 1.667099546E9, 1.667099594E9, 1.667099642E9, 1.66709969E9, 1.667099738E9, 1.667099786E9, 1.667099834E9, 1.667099882E9, 1.66709993E9, 1.667099978E9, 1.667100026E9, 1.667100074E9, 1.667100122E9, 1.66710017E9, 1.667100218E9, 1.667100266E9, 1.667100314E9, 1.667100362E9, 1.66710041E9, 1.667100458E9, 1.667100506E9, 1.667100554E9, 1.667100602E9, 1.66710065E9, 1.66710096E9, 1.66710114E9, 1.667106857E9, 1.667106905E9, 1.667106953E9, 1.667107001E9, 1.667107049E9, 1.667107097E9, 1.667107145E9, 1.667107193E9, 1.667107241E9, 1.667107289E9, 1.667107337E9, 1.667107385E9, 1.667107433E9, 1.667107481E9, 1.667107529E9, 1.667107577E9, 1.667107625E9, 1.667107673E9, 1.667107721E9, 1.667107769E9, 1.667107817E9, 1.667107865E9, 1.667107913E9, 1.667107961E9, 1.667108009E9, 1.667108057E9, 1.667108105E9, 1.667108153E9, 1.667108201E9, 1.667108249E9, 1.667108297E9, 1.667108345E9, 1.667108393E9, 1.667108441E9, 1.667108489E9, 1.667108537E9, 1.667108585E9, 1.667108633E9, 1.667108681E9, 1.667108729E9, 1.667108777E9, 1.667108825E9, 1.667108873E9, 1.667108921E9, 1.667108969E9, 1.667109017E9, 1.667109065E9, 1.667109113E9, 1.667109161E9, 1.667109209E9, 1.667109257E9, 1.667109305E9, 1.667109353E9, 1.667109401E9, 1.667109449E9, 1.667109497E9, 1.667109545E9, 1.667109593E9, 1.667109641E9, 1.667109689E9, 1.667109737E9, 1.667109785E9, 1.667109833E9, 1.667109881E9, 1.667109929E9, 1.667109977E9, 1.667110025E9, 1.667110073E9, 1.667110121E9, 1.667110169E9, 1.6671105E9, 1.66711068E9, 1.667116457E9, 1.667116505E9, 1.667116553E9, 1.667116601E9, 1.667116649E9, 1.667116697E9, 1.667116745E9, 1.667116793E9, 1.667116841E9, 1.667116889E9, 1.667116937E9, 1.667116985E9, 1.667117033E9, 1.667117081E9, 1.667117129E9, 1.667117177E9, 1.667117225E9, 1.667117273E9, 1.667117321E9, 1.667117369E9, 1.667117417E9, 1.667117465E9, 1.667117513E9, 1.667117561E9, 1.667117609E9, 1.667117657E9, 1.667117705E9, 1.667117753E9, 1.667117801E9, 1.667117849E9, 1.667117897E9, 1.667117945E9, 1.667117993E9, 1.667118041E9, 1.667118089E9, 1.667118137E9, 1.667118185E9, 1.667118233E9, 1.667118281E9, 1.667118329E9, 1.667118377E9, 1.667118425E9, 1.667118473E9, 1.667118521E9, 1.667118569E9, 1.667118617E9, 1.667118665E9, 1.667118713E9, 1.667118761E9, 1.667118809E9, 1.667118857E9, 1.667118905E9, 1.667118953E9, 1.667119001E9, 1.667119049E9, 1.667119097E9, 1.667119145E9, 1.667119193E9, 1.667119241E9, 1.667119289E9, 1.667119337E9, 1.667119385E9, 1.667119433E9, 1.667119481E9, 1.667119529E9, 1.6671198E9, 1.66711998E9, 1.667125544E9, 1.667125592E9, 1.66712564E9, 1.667125688E9, 1.667125736E9, 1.667125784E9, 1.667125832E9, 1.66712588E9, 1.667125928E9, 1.667125976E9, 1.667126024E9, 1.667126072E9, 1.66712612E9, 1.667126168E9, 1.667126216E9, 1.667126264E9, 1.667126312E9, 1.66712636E9, 1.667126408E9, 1.667126456E9, 1.667126504E9, 1.667126552E9, 1.6671266E9, 1.667126648E9, 1.667126696E9, 1.667126744E9, 1.667126792E9, 1.66712684E9, 1.667126888E9, 1.667126936E9, 1.667126984E9, 1.667127032E9, 1.66712708E9, 1.667127128E9, 1.667127176E9, 1.667127224E9, 1.667127272E9, 1.66712732E9, 1.667127368E9, 1.667127416E9, 1.667127464E9, 1.667127512E9, 1.66712756E9, 1.667127608E9, 1.667127656E9, 1.667127704E9, 1.667127752E9, 1.6671278E9, 1.667127848E9, 1.667127896E9, 1.667127944E9, 1.667127992E9, 1.66712804E9, 1.667128088E9, 1.667128136E9, 1.667128184E9, 1.667128232E9, 1.66712828E9, 1.667128328E9, 1.667128376E9, 1.667128424E9, 1.667128472E9, 1.66712852E9, 1.667128568E9, 1.667128616E9, 1.667128664E9, 1.667128712E9, 1.66712876E9, 1.6671291E9, 1.66712928E9, 1.667134992E9, 1.66713504E9, 1.667135088E9, 1.667135136E9, 1.667135184E9, 1.667135232E9, 1.66713528E9, 1.667135328E9, 1.667135376E9, 1.667135424E9, 1.667135472E9, 1.66713552E9, 1.667135568E9, 1.667135616E9, 1.667135664E9, 1.667135712E9, 1.66713576E9, 1.667135808E9, 1.667135856E9, 1.667135904E9, 1.667135952E9, 1.667136E9, 1.667136048E9, 1.667136096E9, 1.667136144E9, 1.667136192E9, 1.66713624E9, 1.667136288E9, 1.667136336E9, 1.667136384E9, 1.667136432E9, 1.66713648E9, 1.667136528E9, 1.667136576E9, 1.667136624E9, 1.667136672E9, 1.66713672E9, 1.667136768E9, 1.667136816E9, 1.667136864E9, 1.667136912E9, 1.66713696E9, 1.667137008E9, 1.667137056E9, 1.667137104E9, 1.667137152E9, 1.6671372E9, 1.667137248E9, 1.667137296E9, 1.667137344E9, 1.667137392E9, 1.66713744E9, 1.667137488E9, 1.667137536E9, 1.667137584E9, 1.667137632E9, 1.66713768E9, 1.667137728E9, 1.667137776E9, 1.667137824E9, 1.667137872E9, 1.66713792E9, 1.667137968E9, 1.667138016E9, 1.667138064E9, 1.667138112E9, 1.66713816E9, 1.667138208E9, 1.667138256E9, 1.667138304E9, 1.667138352E9, 1.6671384E9, 1.66713876E9, 1.66713906E9, 1.667144845E9, 1.667144893E9, 1.667144941E9, 1.667144989E9, 1.667145037E9, 1.667145085E9, 1.667145133E9, 1.667145181E9, 1.667145229E9, 1.667145277E9, 1.667145325E9, 1.667145373E9, 1.667145421E9, 1.667145469E9, 1.667145517E9, 1.667145565E9, 1.667145613E9, 1.667145661E9, 1.667145709E9, 1.667145757E9, 1.667145805E9, 1.667145853E9, 1.667145901E9, 1.667145949E9, 1.667145997E9, 1.667146045E9, 1.667146093E9, 1.667146141E9, 1.667146189E9, 1.667146237E9, 1.667146285E9, 1.667146333E9, 1.667146381E9, 1.667146429E9, 1.667146477E9, 1.667146525E9, 1.667146573E9, 1.667146621E9, 1.667146669E9, 1.667146717E9, 1.667146765E9, 1.667146813E9, 1.667146861E9, 1.667146909E9, 1.667146957E9, 1.667147005E9, 1.667147053E9, 1.667147101E9, 1.667147149E9, 1.667147197E9, 1.667147245E9, 1.667147293E9, 1.667147341E9, 1.667147389E9, 1.667147437E9, 1.667147485E9, 1.667147533E9, 1.667147581E9, 1.667147629E9, 1.667147677E9, 1.667147725E9, 1.667147773E9, 1.667147821E9, 1.667147869E9, 1.667147917E9, 1.667147965E9, 1.667148013E9, 1.667148061E9, 1.667148109E9, 1.66714842E9, 1.6671486E9, 1.667154155E9, 1.667154203E9, 1.667154251E9, 1.667154299E9, 1.667154347E9, 1.667154395E9, 1.667154443E9, 1.667154491E9, 1.667154539E9, 1.667154587E9, 1.667154635E9, 1.667154683E9, 1.667154731E9, 1.667154779E9, 1.667154827E9, 1.667154875E9, 1.667154923E9, 1.667154971E9, 1.667155019E9, 1.667155067E9, 1.667155115E9, 1.667155163E9, 1.667155211E9, 1.667155259E9, 1.667155307E9, 1.667155355E9, 1.667155403E9, 1.667155451E9, 1.667155499E9, 1.667155547E9, 1.667155595E9, 1.667155643E9, 1.667155691E9, 1.667155739E9, 1.667155787E9, 1.667155835E9, 1.667155883E9, 1.667155931E9, 1.667155979E9, 1.667156027E9, 1.667156075E9, 1.667156123E9, 1.667156171E9, 1.667156219E9, 1.667156267E9, 1.667156315E9, 1.667156363E9, 1.667156411E9, 1.667156459E9, 1.667156507E9, 1.667156555E9, 1.667156603E9, 1.667156651E9, 1.667156699E9, 1.667156747E9, 1.667156795E9, 1.667156843E9, 1.667156891E9, 1.667156939E9, 1.667156987E9, 1.667157035E9, 1.667157083E9, 1.667157131E9, 1.667157179E9, 1.667157227E9, 1.667157275E9, 1.667157323E9, 1.667157371E9, 1.667157419E9, 1.66715772E9, 1.6671579E9, 1.667163741E9, 1.667163789E9, 1.667163837E9, 1.667163885E9, 1.667163933E9, 1.667163981E9, 1.667164029E9, 1.667164077E9, 1.667164125E9, 1.667164173E9, 1.667164221E9, 1.667164269E9, 1.667164317E9, 1.667164365E9, 1.667164413E9, 1.667164461E9, 1.667164509E9, 1.667164557E9, 1.667164605E9, 1.667164653E9, 1.667164701E9, 1.667164749E9, 1.667164797E9, 1.667164845E9, 1.667164893E9, 1.667164941E9, 1.667164989E9, 1.667165037E9, 1.667165085E9, 1.667165133E9, 1.667165181E9, 1.667165229E9, 1.667165277E9, 1.667165325E9, 1.667165373E9, 1.667165421E9, 1.667165469E9, 1.667165517E9, 1.667165565E9, 1.667165613E9, 1.667165661E9, 1.667165709E9, 1.667165757E9, 1.667165805E9, 1.667165853E9, 1.667165901E9, 1.667165949E9, 1.667165997E9, 1.667166045E9, 1.667166093E9, 1.667166141E9, 1.667166189E9, 1.667166237E9, 1.667166285E9, 1.667166333E9, 1.667166381E9, 1.667166429E9, 1.667166477E9, 1.667166525E9, 1.667166573E9, 1.667166621E9, 1.667166669E9, 1.667166717E9, 1.667166765E9, 1.667166813E9, 1.667166861E9, 1.667166909E9, 1.667166957E9, 1.667167005E9, 1.667167053E9, 1.667167101E9, 1.667167149E9, 1.6671675E9, 1.66716768E9, 1.66717351E9, 1.667173558E9, 1.667173606E9, 1.667173654E9, 1.667173702E9, 1.66717375E9, 1.667173798E9, 1.667173846E9, 1.667173894E9, 1.667173942E9, 1.66717399E9, 1.667174038E9, 1.667174086E9, 1.667174134E9, 1.667174182E9, 1.66717423E9, 1.667174278E9, 1.667174326E9, 1.667174374E9, 1.667174422E9, 1.66717447E9, 1.667174518E9, 1.667174566E9, 1.667174614E9, 1.667174662E9, 1.66717471E9, 1.667174758E9, 1.667174806E9, 1.667174854E9, 1.667174902E9, 1.66717495E9, 1.667174998E9, 1.667175046E9, 1.667175094E9, 1.667175142E9, 1.66717519E9, 1.667175238E9, 1.667175286E9, 1.667175334E9, 1.667175382E9, 1.66717543E9, 1.667175478E9, 1.667175526E9, 1.667175574E9, 1.667175622E9, 1.66717567E9, 1.667175718E9, 1.667175766E9, 1.667175814E9, 1.667175862E9, 1.66717591E9, 1.667175958E9, 1.667176006E9, 1.667176054E9, 1.667176102E9, 1.66717615E9, 1.667176198E9, 1.667176246E9, 1.667176294E9, 1.667176342E9, 1.66717639E9, 1.667176438E9, 1.667176486E9, 1.667176534E9, 1.667176582E9, 1.66717663E9, 1.66717692E9, 1.6671771E9, 1.667182933E9, 1.667182981E9, 1.667183029E9, 1.667183077E9, 1.667183125E9, 1.667183173E9, 1.667183221E9, 1.667183269E9, 1.667183317E9, 1.667183365E9, 1.667183413E9, 1.667183461E9, 1.667183509E9, 1.667183557E9, 1.667183605E9, 1.667183653E9, 1.667183701E9, 1.667183749E9, 1.667183797E9, 1.667183845E9, 1.667183893E9, 1.667183941E9, 1.667183989E9, 1.667184037E9, 1.667184085E9, 1.667184133E9, 1.667184181E9, 1.667184229E9, 1.667184277E9, 1.667184325E9, 1.667184373E9, 1.667184421E9, 1.667184469E9, 1.667184517E9, 1.667184565E9, 1.667184613E9, 1.667184661E9, 1.667184709E9, 1.667184757E9, 1.667184805E9, 1.667184853E9, 1.667184901E9, 1.667184949E9, 1.667184997E9, 1.667185045E9, 1.667185093E9, 1.667185141E9, 1.667185189E9, 1.667185237E9, 1.667185285E9, 1.667185333E9, 1.667185381E9, 1.667185429E9, 1.667185477E9, 1.667185525E9, 1.667185573E9, 1.667185621E9, 1.667185669E9, 1.667185717E9, 1.667185765E9, 1.667185813E9, 1.667185861E9, 1.667185909E9, 1.667185957E9, 1.667186005E9, 1.667186053E9, 1.667186101E9, 1.667186149E9, 1.66718646E9, 1.66718664E9, 1.667192466E9, 1.667192514E9, 1.667192562E9, 1.66719261E9, 1.667192658E9, 1.667192706E9, 1.667192754E9, 1.667192802E9, 1.66719285E9, 1.667192898E9, 1.667192946E9, 1.667192994E9, 1.667193042E9, 1.66719309E9, 1.667193138E9, 1.667193186E9, 1.667193234E9, 1.667193282E9, 1.66719333E9, 1.667193378E9, 1.667193426E9, 1.667193474E9, 1.667193522E9, 1.66719357E9, 1.667193618E9, 1.667193666E9, 1.667193714E9, 1.667193762E9, 1.66719381E9, 1.667193858E9, 1.667193906E9, 1.667193954E9, 1.667194002E9, 1.66719405E9, 1.667194098E9, 1.667194146E9, 1.667194194E9, 1.667194242E9, 1.66719429E9, 1.667194338E9, 1.667194386E9, 1.667194434E9, 1.667194482E9, 1.66719453E9, 1.667194578E9, 1.667194626E9, 1.667194674E9, 1.667194722E9, 1.66719477E9, 1.667194818E9, 1.667194866E9, 1.667194914E9, 1.667194962E9, 1.66719501E9, 1.667195058E9, 1.667195106E9, 1.667195154E9, 1.667195202E9, 1.66719525E9, 1.667195298E9, 1.667195346E9, 1.667195394E9, 1.667195442E9, 1.66719549E9, 1.667195538E9, 1.667195586E9, 1.667195634E9, 1.667195682E9, 1.66719573E9, 1.66719612E9, 1.6671963E9, 1.667202045E9, 1.667202093E9, 1.667202141E9, 1.667202189E9, 1.667202237E9, 1.667202285E9, 1.667202333E9, 1.667202381E9, 1.667202429E9, 1.667202477E9, 1.667202525E9, 1.667202573E9, 1.667202621E9, 1.667202669E9, 1.667202717E9, 1.667202765E9, 1.667202813E9, 1.667202861E9, 1.667202909E9, 1.667202957E9, 1.667203005E9, 1.667203053E9, 1.667203101E9, 1.667203149E9, 1.667203197E9, 1.667203245E9, 1.667203293E9, 1.667203341E9, 1.667203389E9, 1.667203437E9, 1.667203485E9, 1.667203533E9, 1.667203581E9, 1.667203629E9, 1.667203677E9, 1.667203725E9, 1.667203773E9, 1.667203821E9, 1.667203869E9, 1.667203917E9, 1.667203965E9, 1.667204013E9, 1.667204061E9, 1.667204109E9, 1.667204157E9, 1.667204205E9, 1.667204253E9, 1.667204301E9, 1.667204349E9, 1.667204397E9, 1.667204445E9, 1.667204493E9, 1.667204541E9, 1.667204589E9, 1.667204637E9, 1.667204685E9, 1.667204733E9, 1.667204781E9, 1.667204829E9, 1.667204877E9, 1.667204925E9, 1.667204973E9, 1.667205021E9, 1.667205069E9, 1.667205117E9, 1.667205165E9, 1.667205213E9, 1.667205261E9, 1.667205309E9, 1.66720566E9, 1.66720584E9, 1.667211783E9, 1.667211831E9, 1.667211879E9, 1.667211927E9, 1.667211975E9, 1.667212023E9, 1.667212071E9, 1.667212119E9, 1.667212167E9, 1.667212215E9, 1.667212263E9, 1.667212311E9, 1.667212359E9, 1.667212407E9, 1.667212455E9, 1.667212503E9, 1.667212551E9, 1.667212599E9, 1.667212647E9, 1.667212695E9, 1.667212743E9, 1.667212791E9, 1.667212839E9, 1.667212887E9, 1.667212935E9, 1.667212983E9, 1.667213031E9, 1.667213079E9, 1.667213127E9, 1.667213175E9, 1.667213223E9, 1.667213271E9, 1.667213319E9, 1.667213367E9, 1.667213415E9, 1.667213463E9, 1.667213511E9, 1.667213559E9, 1.667213607E9, 1.667213655E9, 1.667213703E9, 1.667213751E9, 1.667213799E9, 1.667213847E9, 1.667213895E9, 1.667213943E9, 1.667213991E9, 1.667214039E9, 1.667214087E9, 1.667214135E9, 1.667214183E9, 1.667214231E9, 1.667214279E9, 1.667214327E9, 1.667214375E9, 1.667214423E9, 1.667214471E9, 1.667214519E9, 1.667214567E9, 1.667214615E9, 1.667214663E9, 1.667214711E9, 1.667214759E9, 1.667214807E9, 1.667214855E9, 1.667214903E9, 1.667214951E9, 1.667214999E9, 1.66721532E9, 1.6672155E9, 1.66722127E9, 1.667221318E9, 1.667221366E9, 1.667221414E9, 1.667221462E9, 1.66722151E9, 1.667221558E9, 1.667221606E9, 1.667221654E9, 1.667221702E9, 1.66722175E9, 1.667221798E9, 1.667221846E9, 1.667221894E9, 1.667221942E9, 1.66722199E9, 1.667222038E9, 1.667222086E9, 1.667222134E9, 1.667222182E9, 1.66722223E9, 1.667222278E9, 1.667222326E9, 1.667222374E9, 1.667222422E9, 1.66722247E9, 1.667222518E9, 1.667222566E9, 1.667222614E9, 1.667222662E9, 1.66722271E9, 1.667222758E9, 1.667222806E9, 1.667222854E9, 1.667222902E9, 1.66722295E9, 1.667222998E9, 1.667223046E9, 1.667223094E9, 1.667223142E9, 1.66722319E9, 1.667223238E9, 1.667223286E9, 1.667223334E9, 1.667223382E9, 1.66722343E9, 1.667223478E9, 1.667223526E9, 1.667223574E9, 1.667223622E9, 1.66722367E9, 1.667223718E9, 1.667223766E9, 1.667223814E9, 1.667223862E9, 1.66722391E9, 1.667223958E9, 1.667224006E9, 1.667224054E9, 1.667224102E9, 1.66722415E9, 1.667224198E9, 1.667224246E9, 1.667224294E9, 1.667224342E9, 1.66722439E9, 1.667224438E9, 1.667224486E9, 1.667224534E9, 1.667224582E9, 1.66722463E9, 1.66722498E9, 1.66722516E9, 1.667231005E9, 1.667231053E9, 1.667231101E9, 1.667231149E9, 1.667231197E9, 1.667231245E9, 1.667231293E9, 1.667231341E9, 1.667231389E9, 1.667231437E9, 1.667231485E9, 1.667231533E9, 1.667231581E9, 1.667231629E9, 1.667231677E9, 1.667231725E9, 1.667231773E9, 1.667231821E9, 1.667231869E9, 1.667231917E9, 1.667231965E9, 1.667232013E9, 1.667232061E9, 1.667232109E9, 1.667232157E9, 1.667232205E9, 1.667232253E9, 1.667232301E9, 1.667232349E9, 1.667232397E9, 1.667232445E9, 1.667232493E9, 1.667232541E9, 1.667232589E9, 1.667232637E9, 1.667232685E9, 1.667232733E9, 1.667232781E9, 1.667232829E9, 1.667232877E9, 1.667232925E9, 1.667232973E9, 1.667233021E9, 1.667233069E9, 1.667233117E9, 1.667233165E9, 1.667233213E9, 1.667233261E9, 1.667233309E9, 1.667233357E9, 1.667233405E9, 1.667233453E9, 1.667233501E9, 1.667233549E9, 1.667233597E9, 1.667233645E9, 1.667233693E9, 1.667233741E9, 1.667233789E9, 1.667233837E9, 1.667233885E9, 1.667233933E9, 1.667233981E9, 1.667234029E9, 1.667234077E9, 1.667234125E9, 1.667234173E9, 1.667234221E9, 1.667234269E9, 1.667234317E9, 1.667234365E9, 1.667234413E9, 1.667234461E9, 1.667234509E9, 1.66723488E9, 1.66723506E9, 1.667240674E9, 1.667240722E9, 1.66724077E9, 1.667240818E9, 1.667240866E9, 1.667240914E9, 1.667240962E9, 1.66724101E9, 1.667241058E9, 1.667241106E9, 1.667241154E9, 1.667241202E9, 1.66724125E9, 1.667241298E9, 1.667241346E9, 1.667241394E9, 1.667241442E9, 1.66724149E9, 1.667241538E9, 1.667241586E9, 1.667241634E9, 1.667241682E9, 1.66724173E9, 1.667241778E9, 1.667241826E9, 1.667241874E9, 1.667241922E9, 1.66724197E9, 1.667242018E9, 1.667242066E9, 1.667242114E9, 1.667242162E9, 1.66724221E9, 1.667242258E9, 1.667242306E9, 1.667242354E9, 1.667242402E9, 1.66724245E9, 1.667242498E9, 1.667242546E9, 1.667242594E9, 1.667242642E9, 1.66724269E9, 1.667242738E9, 1.667242786E9, 1.667242834E9, 1.667242882E9, 1.66724293E9, 1.667242978E9, 1.667243026E9, 1.667243074E9, 1.667243122E9, 1.66724317E9, 1.667243218E9, 1.667243266E9, 1.667243314E9, 1.667243362E9, 1.66724341E9, 1.667243458E9, 1.667243506E9, 1.667243554E9, 1.667243602E9, 1.66724365E9, 1.667243698E9, 1.667243746E9, 1.667243794E9, 1.667243842E9, 1.66724389E9, 1.66724424E9, 1.66724442E9, 1.667250171E9, 1.667250219E9, 1.667250267E9, 1.667250315E9, 1.667250363E9, 1.667250411E9, 1.667250459E9, 1.667250507E9, 1.667250555E9, 1.667250603E9, 1.667250651E9, 1.667250699E9, 1.667250747E9, 1.667250795E9, 1.667250843E9, 1.667250891E9, 1.667250939E9, 1.667250987E9, 1.667251035E9, 1.667251083E9, 1.667251131E9, 1.667251179E9, 1.667251227E9, 1.667251275E9, 1.667251323E9, 1.667251371E9, 1.667251419E9, 1.667251467E9, 1.667251515E9, 1.667251563E9, 1.667251611E9, 1.667251659E9, 1.667251707E9, 1.667251755E9, 1.667251803E9, 1.667251851E9, 1.667251899E9, 1.667251947E9, 1.667251995E9, 1.667252043E9, 1.667252091E9, 1.667252139E9, 1.667252187E9, 1.667252235E9, 1.667252283E9, 1.667252331E9, 1.667252379E9, 1.667252427E9, 1.667252475E9, 1.667252523E9, 1.667252571E9, 1.667252619E9, 1.667252667E9, 1.667252715E9, 1.667252763E9, 1.667252811E9, 1.667252859E9, 1.667252907E9, 1.667252955E9, 1.667253003E9, 1.667253051E9, 1.667253099E9, 1.667253147E9, 1.667253195E9, 1.667253243E9, 1.667253291E9, 1.667253339E9, 1.6672536E9, 1.6672539E9, 1.667259686E9, 1.667259734E9, 1.667259782E9, 1.66725983E9, 1.667259878E9, 1.667259926E9, 1.667259974E9, 1.667260022E9, 1.66726007E9, 1.667260118E9, 1.667260166E9, 1.667260214E9, 1.667260262E9, 1.66726031E9, 1.667260358E9, 1.667260406E9, 1.667260454E9, 1.667260502E9, 1.66726055E9, 1.667260598E9, 1.667260646E9, 1.667260694E9, 1.667260742E9, 1.66726079E9, 1.667260838E9, 1.667260886E9, 1.667260934E9, 1.667260982E9, 1.66726103E9, 1.667261078E9, 1.667261126E9, 1.667261174E9, 1.667261222E9, 1.66726127E9, 1.667261318E9, 1.667261366E9, 1.667261414E9, 1.667261462E9, 1.66726151E9, 1.667261558E9, 1.667261606E9, 1.667261654E9, 1.667261702E9, 1.66726175E9, 1.667261798E9, 1.667261846E9, 1.667261894E9, 1.667261942E9, 1.66726199E9, 1.667262038E9, 1.667262086E9, 1.667262134E9, 1.667262182E9, 1.66726223E9, 1.667262278E9, 1.667262326E9, 1.667262374E9, 1.667262422E9, 1.66726247E9, 1.667262518E9, 1.667262566E9, 1.667262614E9, 1.667262662E9, 1.66726271E9, 1.667262758E9, 1.667262806E9, 1.667262854E9, 1.667262902E9, 1.66726295E9, 1.66726326E9, 1.66726344E9, 1.667269212E9, 1.66726926E9, 1.667269308E9, 1.667269356E9, 1.667269404E9, 1.667269452E9, 1.6672695E9, 1.667269548E9, 1.667269596E9, 1.667269644E9, 1.667269692E9, 1.66726974E9, 1.667269788E9, 1.667269836E9, 1.667269884E9, 1.667269932E9, 1.66726998E9, 1.667270028E9, 1.667270076E9, 1.667270124E9, 1.667270172E9, 1.66727022E9, 1.667270268E9, 1.667270316E9, 1.667270364E9, 1.667270412E9, 1.66727046E9, 1.667270508E9, 1.667270556E9, 1.667270604E9, 1.667270652E9, 1.6672707E9, 1.667270748E9, 1.667270796E9, 1.667270844E9, 1.667270892E9, 1.66727094E9, 1.667270988E9, 1.667271036E9, 1.667271084E9, 1.667271132E9, 1.66727118E9, 1.667271228E9, 1.667271276E9, 1.667271324E9, 1.667271372E9, 1.66727142E9, 1.667271468E9, 1.667271516E9, 1.667271564E9, 1.667271612E9, 1.66727166E9, 1.667271708E9, 1.667271756E9, 1.667271804E9, 1.667271852E9, 1.6672719E9, 1.667271948E9, 1.667271996E9, 1.667272044E9, 1.667272092E9, 1.66727214E9, 1.667272188E9, 1.667272236E9, 1.667272284E9, 1.667272332E9, 1.66727238E9, 1.667272428E9, 1.667272476E9, 1.667272524E9, 1.667272572E9, 1.66727262E9, 1.66727292E9, 1.6672731E9, 1.667278872E9, 1.66727892E9, 1.667278968E9, 1.667279016E9, 1.667279064E9, 1.667279112E9, 1.66727916E9, 1.667279208E9, 1.667279256E9, 1.667279304E9, 1.667279352E9, 1.6672794E9, 1.667279448E9, 1.667279496E9, 1.667279544E9, 1.667279592E9, 1.66727964E9, 1.667279688E9, 1.667279736E9, 1.667279784E9, 1.667279832E9, 1.66727988E9, 1.667279928E9, 1.667279976E9, 1.667280024E9, 1.667280072E9, 1.66728012E9, 1.667280168E9, 1.667280216E9, 1.667280264E9, 1.667280312E9, 1.66728036E9, 1.667280408E9, 1.667280456E9, 1.667280504E9, 1.667280552E9, 1.6672806E9, 1.667280648E9, 1.667280696E9, 1.667280744E9, 1.667280792E9, 1.66728084E9, 1.667280888E9, 1.667280936E9, 1.667280984E9, 1.667281032E9, 1.66728108E9, 1.667281128E9, 1.667281176E9, 1.667281224E9, 1.667281272E9, 1.66728132E9, 1.667281368E9, 1.667281416E9, 1.667281464E9, 1.667281512E9, 1.66728156E9, 1.667281608E9, 1.667281656E9, 1.667281704E9, 1.667281752E9, 1.6672818E9, 1.667281848E9, 1.667281896E9, 1.667281944E9, 1.667281992E9, 1.66728204E9, 1.66728234E9, 1.66728252E9, 1.667288574E9, 1.667288622E9, 1.66728867E9, 1.667288718E9, 1.667288766E9, 1.667288814E9, 1.667288862E9, 1.66728891E9, 1.667288958E9, 1.667289006E9, 1.667289054E9, 1.667289102E9, 1.66728915E9, 1.667289198E9, 1.667289246E9, 1.667289294E9, 1.667289342E9, 1.66728939E9, 1.667289438E9, 1.667289486E9, 1.667289534E9, 1.667289582E9, 1.66728963E9, 1.667289678E9, 1.667289726E9, 1.667289774E9, 1.667289822E9, 1.66728987E9, 1.667289918E9, 1.667289966E9, 1.667290014E9, 1.667290062E9, 1.66729011E9, 1.667290158E9, 1.667290206E9, 1.667290254E9, 1.667290302E9, 1.66729035E9, 1.667290398E9, 1.667290446E9, 1.667290494E9, 1.667290542E9, 1.66729059E9, 1.667290638E9, 1.667290686E9, 1.667290734E9, 1.667290782E9, 1.66729083E9, 1.667290878E9, 1.667290926E9, 1.667290974E9, 1.667291022E9, 1.66729107E9, 1.667291118E9, 1.667291166E9, 1.667291214E9, 1.667291262E9, 1.66729131E9, 1.667291358E9, 1.667291406E9, 1.667291454E9, 1.667291502E9, 1.66729155E9, 1.667291598E9, 1.667291646E9, 1.667291694E9, 1.667291742E9, 1.66729179E9, 1.66729212E9, 1.6672923E9, 1.667298051E9, 1.667298099E9, 1.667298147E9, 1.667298195E9, 1.667298243E9, 1.667298291E9, 1.667298339E9, 1.667298387E9, 1.667298435E9, 1.667298483E9, 1.667298531E9, 1.667298579E9, 1.667298627E9, 1.667298675E9, 1.667298723E9, 1.667298771E9, 1.667298819E9, 1.667298867E9, 1.667298915E9, 1.667298963E9, 1.667299011E9, 1.667299059E9, 1.667299107E9, 1.667299155E9, 1.667299203E9, 1.667299251E9, 1.667299299E9, 1.667299347E9, 1.667299395E9, 1.667299443E9, 1.667299491E9, 1.667299539E9, 1.667299587E9, 1.667299635E9, 1.667299683E9, 1.667299731E9, 1.667299779E9, 1.667299827E9, 1.667299875E9, 1.667299923E9, 1.667299971E9, 1.667300019E9, 1.667300067E9, 1.667300115E9, 1.667300163E9, 1.667300211E9, 1.667300259E9, 1.667300307E9, 1.667300355E9, 1.667300403E9, 1.667300451E9, 1.667300499E9, 1.667300547E9, 1.667300595E9, 1.667300643E9, 1.667300691E9, 1.667300739E9, 1.667300787E9, 1.667300835E9, 1.667300883E9, 1.667300931E9, 1.667300979E9, 1.667301027E9, 1.667301075E9, 1.667301123E9, 1.667301171E9, 1.667301219E9, 1.66730148E9, 1.66730172E9, 1.667307537E9, 1.667307585E9, 1.667307633E9, 1.667307681E9, 1.667307729E9, 1.667307777E9, 1.667307825E9, 1.667307873E9, 1.667307921E9, 1.667307969E9, 1.667308017E9, 1.667308065E9, 1.667308113E9, 1.667308161E9, 1.667308209E9, 1.667308257E9, 1.667308305E9, 1.667308353E9, 1.667308401E9, 1.667308449E9, 1.667308497E9, 1.667308545E9, 1.667308593E9, 1.667308641E9, 1.667308689E9, 1.667308737E9, 1.667308785E9, 1.667308833E9, 1.667308881E9, 1.667308929E9, 1.667308977E9, 1.667309025E9, 1.667309073E9, 1.667309121E9, 1.667309169E9, 1.667309217E9, 1.667309265E9, 1.667309313E9, 1.667309361E9, 1.667309409E9, 1.667309457E9, 1.667309505E9, 1.667309553E9, 1.667309601E9, 1.667309649E9, 1.667309697E9, 1.667309745E9, 1.667309793E9, 1.667309841E9, 1.667309889E9, 1.667309937E9, 1.667309985E9, 1.667310033E9, 1.667310081E9, 1.667310129E9, 1.667310177E9, 1.667310225E9, 1.667310273E9, 1.667310321E9, 1.667310369E9, 1.667310417E9, 1.667310465E9, 1.667310513E9, 1.667310561E9, 1.667310609E9, 1.667310657E9, 1.667310705E9, 1.667310753E9, 1.667310801E9, 1.667310849E9, 1.66731114E9, 1.66731132E9, 1.667317123E9, 1.667317171E9, 1.667317219E9, 1.667317267E9, 1.667317315E9, 1.667317363E9, 1.667317411E9, 1.667317459E9, 1.667317507E9, 1.667317555E9, 1.667317603E9, 1.667317651E9, 1.667317699E9, 1.667317747E9, 1.667317795E9, 1.667317843E9, 1.667317891E9, 1.667317939E9, 1.667317987E9, 1.667318035E9, 1.667318083E9, 1.667318131E9, 1.667318179E9, 1.667318227E9, 1.667318275E9, 1.667318323E9, 1.667318371E9, 1.667318419E9, 1.667318467E9, 1.667318515E9, 1.667318563E9, 1.667318611E9, 1.667318659E9, 1.667318707E9, 1.667318755E9, 1.667318803E9, 1.667318851E9, 1.667318899E9, 1.667318947E9, 1.667318995E9, 1.667319043E9, 1.667319091E9, 1.667319139E9, 1.667319187E9, 1.667319235E9, 1.667319283E9, 1.667319331E9, 1.667319379E9, 1.667319427E9, 1.667319475E9, 1.667319523E9, 1.667319571E9, 1.667319619E9, 1.667319667E9, 1.667319715E9, 1.667319763E9, 1.667319811E9, 1.667319859E9, 1.667319907E9, 1.667319955E9, 1.667320003E9, 1.667320051E9, 1.667320099E9, 1.667320147E9, 1.667320195E9, 1.667320243E9, 1.667320291E9, 1.667320339E9, 1.66732074E9, 1.66732092E9, 1.667326561E9, 1.667326609E9, 1.667326657E9, 1.667326705E9, 1.667326753E9, 1.667326801E9, 1.667326849E9, 1.667326897E9, 1.667326945E9, 1.667326993E9, 1.667327041E9, 1.667327089E9, 1.667327137E9, 1.667327185E9, 1.667327233E9, 1.667327281E9, 1.667327329E9, 1.667327377E9, 1.667327425E9, 1.667327473E9, 1.667327521E9, 1.667327569E9, 1.667327617E9, 1.667327665E9, 1.667327713E9, 1.667327761E9, 1.667327809E9, 1.667327857E9, 1.667327905E9, 1.667327953E9, 1.667328001E9, 1.667328049E9, 1.667328097E9, 1.667328145E9, 1.667328193E9, 1.667328241E9, 1.667328289E9, 1.667328337E9, 1.667328385E9, 1.667328433E9, 1.667328481E9, 1.667328529E9, 1.667328577E9, 1.667328625E9, 1.667328673E9, 1.667328721E9, 1.667328769E9, 1.667328817E9, 1.667328865E9, 1.667328913E9, 1.667328961E9, 1.667329009E9, 1.667329057E9, 1.667329105E9, 1.667329153E9, 1.667329201E9, 1.667329249E9, 1.667329297E9, 1.667329345E9, 1.667329393E9, 1.667329441E9, 1.667329489E9, 1.667329537E9, 1.667329585E9, 1.667329633E9, 1.667329681E9, 1.667329729E9, 1.66733004E9, 1.66733022E9, 1.667335772E9, 1.66733582E9, 1.667335868E9, 1.667335916E9, 1.667335964E9, 1.667336012E9, 1.66733606E9, 1.667336108E9, 1.667336156E9, 1.667336204E9, 1.667336252E9, 1.6673363E9, 1.667336348E9, 1.667336396E9, 1.667336444E9, 1.667336492E9, 1.66733654E9, 1.667336588E9, 1.667336636E9, 1.667336684E9, 1.667336732E9, 1.66733678E9, 1.667336828E9, 1.667336876E9, 1.667336924E9, 1.667336972E9, 1.66733702E9, 1.667337068E9, 1.667337116E9, 1.667337164E9, 1.667337212E9, 1.66733726E9, 1.667337308E9, 1.667337356E9, 1.667337404E9, 1.667337452E9, 1.6673375E9, 1.667337548E9, 1.667337596E9, 1.667337644E9, 1.667337692E9, 1.66733774E9, 1.667337788E9, 1.667337836E9, 1.667337884E9, 1.667337932E9, 1.66733798E9, 1.667338028E9, 1.667338076E9, 1.667338124E9, 1.667338172E9, 1.66733822E9, 1.667338268E9, 1.667338316E9, 1.667338364E9, 1.667338412E9, 1.66733846E9, 1.667338508E9, 1.667338556E9, 1.667338604E9, 1.667338652E9, 1.6673387E9, 1.667338748E9, 1.667338796E9, 1.667338844E9, 1.667338892E9, 1.66733894E9, 1.667338988E9, 1.667339036E9, 1.667339084E9, 1.667339132E9, 1.66733918E9, 1.66733958E9, 1.66733976E9, 1.667345516E9, 1.667345564E9, 1.667345612E9, 1.66734566E9, 1.667345708E9, 1.667345756E9, 1.667345804E9, 1.667345852E9, 1.6673459E9, 1.667345948E9, 1.667345996E9, 1.667346044E9, 1.667346092E9, 1.66734614E9, 1.667346188E9, 1.667346236E9, 1.667346284E9, 1.667346332E9, 1.66734638E9, 1.667346428E9, 1.667346476E9, 1.667346524E9, 1.667346572E9, 1.66734662E9, 1.667346668E9, 1.667346716E9, 1.667346764E9, 1.667346812E9, 1.66734686E9, 1.667346908E9, 1.667346956E9, 1.667347004E9, 1.667347052E9, 1.6673471E9, 1.667347148E9, 1.667347196E9, 1.667347244E9, 1.667347292E9, 1.66734734E9, 1.667347388E9, 1.667347436E9, 1.667347484E9, 1.667347532E9, 1.66734758E9, 1.667347628E9, 1.667347676E9, 1.667347724E9, 1.667347772E9, 1.66734782E9, 1.667347868E9, 1.667347916E9, 1.667347964E9, 1.667348012E9, 1.66734806E9, 1.667348108E9, 1.667348156E9, 1.667348204E9, 1.667348252E9, 1.6673483E9, 1.667348348E9, 1.667348396E9, 1.667348444E9, 1.667348492E9, 1.66734854E9, 1.667348588E9, 1.667348636E9, 1.667348684E9, 1.667348732E9, 1.66734878E9, 1.66734918E9, 1.667349181E9, 1.667354913E9, 1.667354961E9, 1.667355009E9, 1.667355057E9, 1.667355105E9, 1.667355153E9, 1.667355201E9, 1.667355249E9, 1.667355297E9, 1.667355345E9, 1.667355393E9, 1.667355441E9, 1.667355489E9, 1.667355537E9, 1.667355585E9, 1.667355633E9, 1.667355681E9, 1.667355729E9, 1.667355777E9, 1.667355825E9, 1.667355873E9, 1.667355921E9, 1.667355969E9, 1.667356017E9, 1.667356065E9, 1.667356113E9, 1.667356161E9, 1.667356209E9, 1.667356257E9, 1.667356305E9, 1.667356353E9, 1.667356401E9, 1.667356449E9, 1.667356497E9, 1.667356545E9, 1.667356593E9, 1.667356641E9, 1.667356689E9, 1.667356737E9, 1.667356785E9, 1.667356833E9, 1.667356881E9, 1.667356929E9, 1.667356977E9, 1.667357025E9, 1.667357073E9, 1.667357121E9, 1.667357169E9, 1.667357217E9, 1.667357265E9, 1.667357313E9, 1.667357361E9, 1.667357409E9, 1.667357457E9, 1.667357505E9, 1.667357553E9, 1.667357601E9, 1.667357649E9, 1.667357697E9, 1.667357745E9, 1.667357793E9, 1.667357841E9, 1.667357889E9, 1.667357937E9, 1.667357985E9, 1.667358033E9, 1.667358081E9, 1.667358129E9, 1.66735842E9, 1.6673586E9, 1.667364289E9, 1.667364337E9, 1.667364385E9, 1.667364433E9, 1.667364481E9, 1.667364529E9, 1.667364577E9, 1.667364625E9, 1.667364673E9, 1.667364721E9, 1.667364769E9, 1.667364817E9, 1.667364865E9, 1.667364913E9, 1.667364961E9, 1.667365009E9, 1.667365057E9, 1.667365105E9, 1.667365153E9, 1.667365201E9, 1.667365249E9, 1.667365297E9, 1.667365345E9, 1.667365393E9, 1.667365441E9, 1.667365489E9, 1.667365537E9, 1.667365585E9, 1.667365633E9, 1.667365681E9, 1.667365729E9, 1.667365777E9, 1.667365825E9, 1.667365873E9, 1.667365921E9, 1.667365969E9, 1.667366017E9, 1.667366065E9, 1.667366113E9, 1.667366161E9, 1.667366209E9, 1.667366257E9, 1.667366305E9, 1.667366353E9, 1.667366401E9, 1.667366449E9, 1.667366497E9, 1.667366545E9, 1.667366593E9, 1.667366641E9, 1.667366689E9, 1.667366737E9, 1.667366785E9, 1.667366833E9, 1.667366881E9, 1.667366929E9, 1.667366977E9, 1.667367025E9, 1.667367073E9, 1.667367121E9, 1.667367169E9, 1.667367217E9, 1.667367265E9, 1.667367313E9, 1.667367361E9, 1.667367409E9, 1.667367457E9, 1.667367505E9, 1.667367553E9, 1.667367601E9, 1.667367649E9, 1.66736796E9, 1.66736814E9, 1.667373703E9, 1.667373751E9, 1.667373799E9, 1.667373847E9, 1.667373895E9, 1.667373943E9, 1.667373991E9, 1.667374039E9, 1.667374087E9, 1.667374135E9, 1.667374183E9, 1.667374231E9, 1.667374279E9, 1.667374327E9, 1.667374375E9, 1.667374423E9, 1.667374471E9, 1.667374519E9, 1.667374567E9, 1.667374615E9, 1.667374663E9, 1.667374711E9, 1.667374759E9, 1.667374807E9, 1.667374855E9, 1.667374903E9, 1.667374951E9, 1.667374999E9, 1.667375047E9, 1.667375095E9, 1.667375143E9, 1.667375191E9, 1.667375239E9, 1.667375287E9, 1.667375335E9, 1.667375383E9, 1.667375431E9, 1.667375479E9, 1.667375527E9, 1.667375575E9, 1.667375623E9, 1.667375671E9, 1.667375719E9, 1.667375767E9, 1.667375815E9, 1.667375863E9, 1.667375911E9, 1.667375959E9, 1.667376007E9, 1.667376055E9, 1.667376103E9, 1.667376151E9, 1.667376199E9, 1.667376247E9, 1.667376295E9, 1.667376343E9, 1.667376391E9, 1.667376439E9, 1.667376487E9, 1.667376535E9, 1.667376583E9, 1.667376631E9, 1.667376679E9, 1.667376727E9, 1.667376775E9, 1.667376823E9, 1.667376871E9, 1.667376919E9, 1.66737732E9, 1.6673775E9, 1.667383184E9, 1.667383232E9, 1.66738328E9, 1.667383328E9, 1.667383376E9, 1.667383424E9, 1.667383472E9, 1.66738352E9, 1.667383568E9, 1.667383616E9, 1.667383664E9, 1.667383712E9, 1.66738376E9, 1.667383808E9, 1.667383856E9, 1.667383904E9, 1.667383952E9, 1.667384E9, 1.667384048E9, 1.667384096E9, 1.667384144E9, 1.667384192E9, 1.66738424E9, 1.667384288E9, 1.667384336E9, 1.667384384E9, 1.667384432E9, 1.66738448E9, 1.667384528E9, 1.667384576E9, 1.667384624E9, 1.667384672E9, 1.66738472E9, 1.667384768E9, 1.667384816E9, 1.667384864E9, 1.667384912E9, 1.66738496E9, 1.667385008E9, 1.667385056E9, 1.667385104E9, 1.667385152E9, 1.6673852E9, 1.667385248E9, 1.667385296E9, 1.667385344E9, 1.667385392E9, 1.66738544E9, 1.667385488E9, 1.667385536E9, 1.667385584E9, 1.667385632E9, 1.66738568E9, 1.667385728E9, 1.667385776E9, 1.667385824E9, 1.667385872E9, 1.66738592E9, 1.667385968E9, 1.667386016E9, 1.667386064E9, 1.667386112E9, 1.66738616E9, 1.667386208E9, 1.667386256E9, 1.667386304E9, 1.667386352E9, 1.6673864E9, 1.66738668E9, 1.66738686E9, 1.667392473E9, 1.667392521E9, 1.667392569E9, 1.667392617E9, 1.667392665E9, 1.667392713E9, 1.667392761E9, 1.667392809E9, 1.667392857E9, 1.667392905E9, 1.667392953E9, 1.667393001E9, 1.667393049E9, 1.667393097E9, 1.667393145E9, 1.667393193E9, 1.667393241E9, 1.667393289E9, 1.667393337E9, 1.667393385E9, 1.667393433E9, 1.667393481E9, 1.667393529E9, 1.667393577E9, 1.667393625E9, 1.667393673E9, 1.667393721E9, 1.667393769E9, 1.667393817E9, 1.667393865E9, 1.667393913E9, 1.667393961E9, 1.667394009E9, 1.667394057E9, 1.667394105E9, 1.667394153E9, 1.667394201E9, 1.667394249E9, 1.667394297E9, 1.667394345E9, 1.667394393E9, 1.667394441E9, 1.667394489E9, 1.667394537E9, 1.667394585E9, 1.667394633E9, 1.667394681E9, 1.667394729E9, 1.667394777E9, 1.667394825E9, 1.667394873E9, 1.667394921E9, 1.667394969E9, 1.667395017E9, 1.667395065E9, 1.667395113E9, 1.667395161E9, 1.667395209E9, 1.667395257E9, 1.667395305E9, 1.667395353E9, 1.667395401E9, 1.667395449E9, 1.667395497E9, 1.667395545E9, 1.667395593E9, 1.667395641E9, 1.667395689E9, 1.667395737E9, 1.667395785E9, 1.667395833E9, 1.667395881E9, 1.667395929E9, 1.66739616E9, 1.66739634E9, 1.6674024E9, 1.667402448E9, 1.667402496E9, 1.667402544E9, 1.667402592E9, 1.66740264E9, 1.667402688E9, 1.667402736E9, 1.667402784E9, 1.667402832E9, 1.66740288E9, 1.667402928E9, 1.667402976E9, 1.667403024E9, 1.667403072E9, 1.66740312E9, 1.667403168E9, 1.667403216E9, 1.667403264E9, 1.667403312E9, 1.66740336E9, 1.667403408E9, 1.667403456E9, 1.667403504E9, 1.667403552E9, 1.6674036E9, 1.667403648E9, 1.667403696E9, 1.667403744E9, 1.667403792E9, 1.66740384E9, 1.667403888E9, 1.667403936E9, 1.667403984E9, 1.667404032E9, 1.66740408E9, 1.667404128E9, 1.667404176E9, 1.667404224E9, 1.667404272E9, 1.66740432E9, 1.667404368E9, 1.667404416E9, 1.667404464E9, 1.667404512E9, 1.66740456E9, 1.667404608E9, 1.667404656E9, 1.667404704E9, 1.667404752E9, 1.6674048E9, 1.667404848E9, 1.667404896E9, 1.667404944E9, 1.667404992E9, 1.66740504E9, 1.667405088E9, 1.667405136E9, 1.667405184E9, 1.667405232E9, 1.66740528E9, 1.667405328E9, 1.667405376E9, 1.667405424E9, 1.667405472E9, 1.66740552E9, 1.66740588E9, 1.667405881E9, 1.667411575E9, 1.667411623E9, 1.667411671E9, 1.667411719E9, 1.667411767E9, 1.667411815E9, 1.667411863E9, 1.667411911E9, 1.667411959E9, 1.667412007E9, 1.667412055E9, 1.667412103E9, 1.667412151E9, 1.667412199E9, 1.667412247E9, 1.667412295E9, 1.667412343E9, 1.667412391E9, 1.667412439E9, 1.667412487E9, 1.667412535E9, 1.667412583E9, 1.667412631E9, 1.667412679E9, 1.667412727E9, 1.667412775E9, 1.667412823E9, 1.667412871E9, 1.667412919E9, 1.667412967E9, 1.667413015E9, 1.667413063E9, 1.667413111E9, 1.667413159E9, 1.667413207E9, 1.667413255E9, 1.667413303E9, 1.667413351E9, 1.667413399E9, 1.667413447E9, 1.667413495E9, 1.667413543E9, 1.667413591E9, 1.667413639E9, 1.667413687E9, 1.667413735E9, 1.667413783E9, 1.667413831E9, 1.667413879E9, 1.667413927E9, 1.667413975E9, 1.667414023E9, 1.667414071E9, 1.667414119E9, 1.667414167E9, 1.667414215E9, 1.667414263E9, 1.667414311E9, 1.667414359E9, 1.667414407E9, 1.667414455E9, 1.667414503E9, 1.667414551E9, 1.667414599E9, 1.667414647E9, 1.667414695E9, 1.667414743E9, 1.667414791E9, 1.667414839E9, 1.66741512E9, 1.6674153E9, 1.667420981E9, 1.667421029E9, 1.667421077E9, 1.667421125E9, 1.667421173E9, 1.667421221E9, 1.667421269E9, 1.667421317E9, 1.667421365E9, 1.667421413E9, 1.667421461E9, 1.667421509E9, 1.667421557E9, 1.667421605E9, 1.667421653E9, 1.667421701E9, 1.667421749E9, 1.667421797E9, 1.667421845E9, 1.667421893E9, 1.667421941E9, 1.667421989E9, 1.667422037E9, 1.667422085E9, 1.667422133E9, 1.667422181E9, 1.667422229E9, 1.667422277E9, 1.667422325E9, 1.667422373E9, 1.667422421E9, 1.667422469E9, 1.667422517E9, 1.667422565E9, 1.667422613E9, 1.667422661E9, 1.667422709E9, 1.667422757E9, 1.667422805E9, 1.667422853E9, 1.667422901E9, 1.667422949E9, 1.667422997E9, 1.667423045E9, 1.667423093E9, 1.667423141E9, 1.667423189E9, 1.667423237E9, 1.667423285E9, 1.667423333E9, 1.667423381E9, 1.667423429E9, 1.667423477E9, 1.667423525E9, 1.667423573E9, 1.667423621E9, 1.667423669E9, 1.667423717E9, 1.667423765E9, 1.667423813E9, 1.667423861E9, 1.667423909E9, 1.667423957E9, 1.667424005E9, 1.667424053E9, 1.667424101E9, 1.667424149E9, 1.667424197E9, 1.667424245E9, 1.667424293E9, 1.667424341E9, 1.667424389E9, 1.66742472E9, 1.6674249E9, 1.667430619E9, 1.667430667E9, 1.667430715E9, 1.667430763E9, 1.667430811E9, 1.667430859E9, 1.667430907E9, 1.667430955E9, 1.667431003E9, 1.667431051E9, 1.667431099E9, 1.667431147E9, 1.667431195E9, 1.667431243E9, 1.667431291E9, 1.667431339E9, 1.667431387E9, 1.667431435E9, 1.667431483E9, 1.667431531E9, 1.667431579E9, 1.667431627E9, 1.667431675E9, 1.667431723E9, 1.667431771E9, 1.667431819E9, 1.667431867E9, 1.667431915E9, 1.667431963E9, 1.667432011E9, 1.667432059E9, 1.667432107E9, 1.667432155E9, 1.667432203E9, 1.667432251E9, 1.667432299E9, 1.667432347E9, 1.667432395E9, 1.667432443E9, 1.667432491E9, 1.667432539E9, 1.667432587E9, 1.667432635E9, 1.667432683E9, 1.667432731E9, 1.667432779E9, 1.667432827E9, 1.667432875E9, 1.667432923E9, 1.667432971E9, 1.667433019E9, 1.667433067E9, 1.667433115E9, 1.667433163E9, 1.667433211E9, 1.667433259E9, 1.667433307E9, 1.667433355E9, 1.667433403E9, 1.667433451E9, 1.667433499E9, 1.667433547E9, 1.667433595E9, 1.667433643E9, 1.667433691E9, 1.667433739E9, 1.667433787E9, 1.667433835E9, 1.667433883E9, 1.667433931E9, 1.667433979E9, 1.66743432E9, 1.6674345E9, 1.667440053E9, 1.667440101E9, 1.667440149E9, 1.667440197E9, 1.667440245E9, 1.667440293E9, 1.667440341E9, 1.667440389E9, 1.667440437E9, 1.667440485E9, 1.667440533E9, 1.667440581E9, 1.667440629E9, 1.667440677E9, 1.667440725E9, 1.667440773E9, 1.667440821E9, 1.667440869E9, 1.667440917E9, 1.667440965E9, 1.667441013E9, 1.667441061E9, 1.667441109E9, 1.667441157E9, 1.667441205E9, 1.667441253E9, 1.667441301E9, 1.667441349E9, 1.667441397E9, 1.667441445E9, 1.667441493E9, 1.667441541E9, 1.667441589E9, 1.667441637E9, 1.667441685E9, 1.667441733E9, 1.667441781E9, 1.667441829E9, 1.667441877E9, 1.667441925E9, 1.667441973E9, 1.667442021E9, 1.667442069E9, 1.667442117E9, 1.667442165E9, 1.667442213E9, 1.667442261E9, 1.667442309E9, 1.667442357E9, 1.667442405E9, 1.667442453E9, 1.667442501E9, 1.667442549E9, 1.667442597E9, 1.667442645E9, 1.667442693E9, 1.667442741E9, 1.667442789E9, 1.667442837E9, 1.667442885E9, 1.667442933E9, 1.667442981E9, 1.667443029E9, 1.667443077E9, 1.667443125E9, 1.667443173E9, 1.667443221E9, 1.667443269E9, 1.667443317E9, 1.667443365E9, 1.667443413E9, 1.667443461E9, 1.667443509E9, 1.66744374E9, 1.66744392E9, 1.667449653E9, 1.667449701E9, 1.667449749E9, 1.667449797E9, 1.667449845E9, 1.667449893E9, 1.667449941E9, 1.667449989E9, 1.667450037E9, 1.667450085E9, 1.667450133E9, 1.667450181E9, 1.667450229E9, 1.667450277E9, 1.667450325E9, 1.667450373E9, 1.667450421E9, 1.667450469E9, 1.667450517E9, 1.667450565E9, 1.667450613E9, 1.667450661E9, 1.667450709E9, 1.667450757E9, 1.667450805E9, 1.667450853E9, 1.667450901E9, 1.667450949E9, 1.667450997E9, 1.667451045E9, 1.667451093E9, 1.667451141E9, 1.667451189E9, 1.667451237E9, 1.667451285E9, 1.667451333E9, 1.667451381E9, 1.667451429E9, 1.667451477E9, 1.667451525E9, 1.667451573E9, 1.667451621E9, 1.667451669E9, 1.667451717E9, 1.667451765E9, 1.667451813E9, 1.667451861E9, 1.667451909E9, 1.667451957E9, 1.667452005E9, 1.667452053E9, 1.667452101E9, 1.667452149E9, 1.667452197E9, 1.667452245E9, 1.667452293E9, 1.667452341E9, 1.667452389E9, 1.667452437E9, 1.667452485E9, 1.667452533E9, 1.667452581E9, 1.667452629E9, 1.667452677E9, 1.667452725E9, 1.667452773E9, 1.667452821E9, 1.667452869E9, 1.667452917E9, 1.667452965E9, 1.667453013E9, 1.667453061E9, 1.667453109E9, 1.6674534E9, 1.66745358E9, 1.667459184E9, 1.667459232E9, 1.66745928E9, 1.667459328E9, 1.667459376E9, 1.667459424E9, 1.667459472E9, 1.66745952E9, 1.667459568E9, 1.667459616E9, 1.667459664E9, 1.667459712E9, 1.66745976E9, 1.667459808E9, 1.667459856E9, 1.667459904E9, 1.667459952E9, 1.66746E9, 1.667460048E9, 1.667460096E9, 1.667460144E9, 1.667460192E9, 1.66746024E9, 1.667460288E9, 1.667460336E9, 1.667460384E9, 1.667460432E9, 1.66746048E9, 1.667460528E9, 1.667460576E9, 1.667460624E9, 1.667460672E9, 1.66746072E9, 1.667460768E9, 1.667460816E9, 1.667460864E9, 1.667460912E9, 1.66746096E9, 1.667461008E9, 1.667461056E9, 1.667461104E9, 1.667461152E9, 1.6674612E9, 1.667461248E9, 1.667461296E9, 1.667461344E9, 1.667461392E9, 1.66746144E9, 1.667461488E9, 1.667461536E9, 1.667461584E9, 1.667461632E9, 1.66746168E9, 1.667461728E9, 1.667461776E9, 1.667461824E9, 1.667461872E9, 1.66746192E9, 1.667461968E9, 1.667462016E9, 1.667462064E9, 1.667462112E9, 1.66746216E9, 1.667462208E9, 1.667462256E9, 1.667462304E9, 1.667462352E9, 1.6674624E9, 1.66746276E9, 1.66746294E9, 1.667468544E9, 1.667468592E9, 1.66746864E9, 1.667468688E9, 1.667468736E9, 1.667468784E9, 1.667468832E9, 1.66746888E9, 1.667468928E9, 1.667468976E9, 1.667469024E9, 1.667469072E9, 1.66746912E9, 1.667469168E9, 1.667469216E9, 1.667469264E9, 1.667469312E9, 1.66746936E9, 1.667469408E9, 1.667469456E9, 1.667469504E9, 1.667469552E9, 1.6674696E9, 1.667469648E9, 1.667469696E9, 1.667469744E9, 1.667469792E9, 1.66746984E9, 1.667469888E9, 1.667469936E9, 1.667469984E9, 1.667470032E9, 1.66747008E9, 1.667470128E9, 1.667470176E9, 1.667470224E9, 1.667470272E9, 1.66747032E9, 1.667470368E9, 1.667470416E9, 1.667470464E9, 1.667470512E9, 1.66747056E9, 1.667470608E9, 1.667470656E9, 1.667470704E9, 1.667470752E9, 1.6674708E9, 1.667470848E9, 1.667470896E9, 1.667470944E9, 1.667470992E9, 1.66747104E9, 1.667471088E9, 1.667471136E9, 1.667471184E9, 1.667471232E9, 1.66747128E9, 1.667471328E9, 1.667471376E9, 1.667471424E9, 1.667471472E9, 1.66747152E9, 1.667471568E9, 1.667471616E9, 1.667471664E9, 1.667471712E9, 1.66747176E9, 1.66747206E9, 1.66747224E9, 1.667477954E9, 1.667478002E9, 1.66747805E9, 1.667478098E9, 1.667478146E9, 1.667478194E9, 1.667478242E9, 1.66747829E9, 1.667478338E9, 1.667478386E9, 1.667478434E9, 1.667478482E9, 1.66747853E9, 1.667478578E9, 1.667478626E9, 1.667478674E9, 1.667478722E9, 1.66747877E9, 1.667478818E9, 1.667478866E9, 1.667478914E9, 1.667478962E9, 1.66747901E9, 1.667479058E9, 1.667479106E9, 1.667479154E9, 1.667479202E9, 1.66747925E9, 1.667479298E9, 1.667479346E9, 1.667479394E9, 1.667479442E9, 1.66747949E9, 1.667479538E9, 1.667479586E9, 1.667479634E9, 1.667479682E9, 1.66747973E9, 1.667479778E9, 1.667479826E9, 1.667479874E9, 1.667479922E9, 1.66747997E9, 1.667480018E9, 1.667480066E9, 1.667480114E9, 1.667480162E9, 1.66748021E9, 1.667480258E9, 1.667480306E9, 1.667480354E9, 1.667480402E9, 1.66748045E9, 1.667480498E9, 1.667480546E9, 1.667480594E9, 1.667480642E9, 1.66748069E9, 1.667480738E9, 1.667480786E9, 1.667480834E9, 1.667480882E9, 1.66748093E9, 1.667480978E9, 1.667481026E9, 1.667481074E9, 1.667481122E9, 1.66748117E9, 1.66748148E9, 1.66748166E9, 1.667487566E9, 1.667487614E9, 1.667487662E9, 1.66748771E9, 1.667487758E9, 1.667487806E9, 1.667487854E9, 1.667487902E9, 1.66748795E9, 1.667487998E9, 1.667488046E9, 1.667488094E9, 1.667488142E9, 1.66748819E9, 1.667488238E9, 1.667488286E9, 1.667488334E9, 1.667488382E9, 1.66748843E9, 1.667488478E9, 1.667488526E9, 1.667488574E9, 1.667488622E9, 1.66748867E9, 1.667488718E9, 1.667488766E9, 1.667488814E9, 1.667488862E9, 1.66748891E9, 1.667488958E9, 1.667489006E9, 1.667489054E9, 1.667489102E9, 1.66748915E9, 1.667489198E9, 1.667489246E9, 1.667489294E9, 1.667489342E9, 1.66748939E9, 1.667489438E9, 1.667489486E9, 1.667489534E9, 1.667489582E9, 1.66748963E9, 1.667489678E9, 1.667489726E9, 1.667489774E9, 1.667489822E9, 1.66748987E9, 1.667489918E9, 1.667489966E9, 1.667490014E9, 1.667490062E9, 1.66749011E9, 1.667490158E9, 1.667490206E9, 1.667490254E9, 1.667490302E9, 1.66749035E9, 1.667490398E9, 1.667490446E9, 1.667490494E9, 1.667490542E9, 1.66749059E9, 1.667490638E9, 1.667490686E9, 1.667490734E9, 1.667490782E9, 1.66749083E9, 1.66749114E9, 1.66749132E9, 1.66749688E9, 1.667496928E9, 1.667496976E9, 1.667497024E9, 1.667497072E9, 1.66749712E9, 1.667497168E9, 1.667497216E9, 1.667497264E9, 1.667497312E9, 1.66749736E9, 1.667497408E9, 1.667497456E9, 1.667497504E9, 1.667497552E9, 1.6674976E9, 1.667497648E9, 1.667497696E9, 1.667497744E9, 1.667497792E9, 1.66749784E9, 1.667497888E9, 1.667497936E9, 1.667497984E9, 1.667498032E9, 1.66749808E9, 1.667498128E9, 1.667498176E9, 1.667498224E9, 1.667498272E9, 1.66749832E9, 1.667498368E9, 1.667498416E9, 1.667498464E9, 1.667498512E9, 1.66749856E9, 1.667498608E9, 1.667498656E9, 1.667498704E9, 1.667498752E9, 1.6674988E9, 1.667498848E9, 1.667498896E9, 1.667498944E9, 1.667498992E9, 1.66749904E9, 1.667499088E9, 1.667499136E9, 1.667499184E9, 1.667499232E9, 1.66749928E9, 1.667499328E9, 1.667499376E9, 1.667499424E9, 1.667499472E9, 1.66749952E9, 1.667499568E9, 1.667499616E9, 1.667499664E9, 1.667499712E9, 1.66749976E9, 1.667499808E9, 1.667499856E9, 1.667499904E9, 1.667499952E9, 1.6675E9, 1.667500048E9, 1.667500096E9, 1.667500144E9, 1.667500192E9, 1.66750024E9, 1.66750056E9, 1.66750074E9, 1.667506564E9, 1.667506612E9, 1.66750666E9, 1.667506708E9, 1.667506756E9, 1.667506804E9, 1.667506852E9, 1.6675069E9, 1.667506948E9, 1.667506996E9, 1.667507044E9, 1.667507092E9, 1.66750714E9, 1.667507188E9, 1.667507236E9, 1.667507284E9, 1.667507332E9, 1.66750738E9, 1.667507428E9, 1.667507476E9, 1.667507524E9, 1.667507572E9, 1.66750762E9, 1.667507668E9, 1.667507716E9, 1.667507764E9, 1.667507812E9, 1.66750786E9, 1.667507908E9, 1.667507956E9, 1.667508004E9, 1.667508052E9, 1.6675081E9, 1.667508148E9, 1.667508196E9, 1.667508244E9, 1.667508292E9, 1.66750834E9, 1.667508388E9, 1.667508436E9, 1.667508484E9, 1.667508532E9, 1.66750858E9, 1.667508628E9, 1.667508676E9, 1.667508724E9, 1.667508772E9, 1.66750882E9, 1.667508868E9, 1.667508916E9, 1.667508964E9, 1.667509012E9, 1.66750906E9, 1.667509108E9, 1.667509156E9, 1.667509204E9, 1.667509252E9, 1.6675093E9, 1.667509348E9, 1.667509396E9, 1.667509444E9, 1.667509492E9, 1.66750954E9, 1.667509588E9, 1.667509636E9, 1.667509684E9, 1.667509732E9, 1.66750978E9, 1.66751016E9, 1.66751028E9, 1.667515867E9, 1.667515915E9, 1.667515963E9, 1.667516011E9, 1.667516059E9, 1.667516107E9, 1.667516155E9, 1.667516203E9, 1.667516251E9, 1.667516299E9, 1.667516347E9, 1.667516395E9, 1.667516443E9, 1.667516491E9, 1.667516539E9, 1.667516587E9, 1.667516635E9, 1.667516683E9, 1.667516731E9, 1.667516779E9, 1.667516827E9, 1.667516875E9, 1.667516923E9, 1.667516971E9, 1.667517019E9, 1.667517067E9, 1.667517115E9, 1.667517163E9, 1.667517211E9, 1.667517259E9, 1.667517307E9, 1.667517355E9, 1.667517403E9, 1.667517451E9, 1.667517499E9, 1.667517547E9, 1.667517595E9, 1.667517643E9, 1.667517691E9, 1.667517739E9, 1.667517787E9, 1.667517835E9, 1.667517883E9, 1.667517931E9, 1.667517979E9, 1.667518027E9, 1.667518075E9, 1.667518123E9, 1.667518171E9, 1.667518219E9, 1.667518267E9, 1.667518315E9, 1.667518363E9, 1.667518411E9, 1.667518459E9, 1.667518507E9, 1.667518555E9, 1.667518603E9, 1.667518651E9, 1.667518699E9, 1.667518747E9, 1.667518795E9, 1.667518843E9, 1.667518891E9, 1.667518939E9, 1.667518987E9, 1.667519035E9, 1.667519083E9, 1.667519131E9, 1.667519179E9, 1.66751952E9, 1.6675197E9, 1.667525152E9, 1.6675252E9, 1.667525248E9, 1.667525296E9, 1.667525344E9, 1.667525392E9, 1.66752544E9, 1.667525488E9, 1.667525536E9, 1.667525584E9, 1.667525632E9, 1.66752568E9, 1.667525728E9, 1.667525776E9, 1.667525824E9, 1.667525872E9, 1.66752592E9, 1.667525968E9, 1.667526016E9, 1.667526064E9, 1.667526112E9, 1.66752616E9, 1.667526208E9, 1.667526256E9, 1.667526304E9, 1.667526352E9, 1.6675264E9, 1.667526448E9, 1.667526496E9, 1.667526544E9, 1.667526592E9, 1.66752664E9, 1.667526688E9, 1.667526736E9, 1.667526784E9, 1.667526832E9, 1.66752688E9, 1.667526928E9, 1.667526976E9, 1.667527024E9, 1.667527072E9, 1.66752712E9, 1.667527168E9, 1.667527216E9, 1.667527264E9, 1.667527312E9, 1.66752736E9, 1.667527408E9, 1.667527456E9, 1.667527504E9, 1.667527552E9, 1.6675276E9, 1.667527648E9, 1.667527696E9, 1.667527744E9, 1.667527792E9, 1.66752784E9, 1.667527888E9, 1.667527936E9, 1.667527984E9, 1.667528032E9, 1.66752808E9, 1.667528128E9, 1.667528176E9, 1.667528224E9, 1.667528272E9, 1.66752832E9, 1.6675287E9, 1.66752894E9, 1.667534647E9, 1.667534695E9, 1.667534743E9, 1.667534791E9, 1.667534839E9, 1.667534887E9, 1.667534935E9, 1.667534983E9, 1.667535031E9, 1.667535079E9, 1.667535127E9, 1.667535175E9, 1.667535223E9, 1.667535271E9, 1.667535319E9, 1.667535367E9, 1.667535415E9, 1.667535463E9, 1.667535511E9, 1.667535559E9, 1.667535607E9, 1.667535655E9, 1.667535703E9, 1.667535751E9, 1.667535799E9, 1.667535847E9, 1.667535895E9, 1.667535943E9, 1.667535991E9, 1.667536039E9, 1.667536087E9, 1.667536135E9, 1.667536183E9, 1.667536231E9, 1.667536279E9, 1.667536327E9, 1.667536375E9, 1.667536423E9, 1.667536471E9, 1.667536519E9, 1.667536567E9, 1.667536615E9, 1.667536663E9, 1.667536711E9, 1.667536759E9, 1.667536807E9, 1.667536855E9, 1.667536903E9, 1.667536951E9, 1.667536999E9, 1.667537047E9, 1.667537095E9, 1.667537143E9, 1.667537191E9, 1.667537239E9, 1.667537287E9, 1.667537335E9, 1.667537383E9, 1.667537431E9, 1.667537479E9, 1.667537527E9, 1.667537575E9, 1.667537623E9, 1.667537671E9, 1.667537719E9, 1.667537767E9, 1.667537815E9, 1.667537863E9, 1.667537911E9, 1.667537959E9, 1.66753824E9, 1.66753842E9, 1.667544105E9, 1.667544153E9, 1.667544201E9, 1.667544249E9, 1.667544297E9, 1.667544345E9, 1.667544393E9, 1.667544441E9, 1.667544489E9, 1.667544537E9, 1.667544585E9, 1.667544633E9, 1.667544681E9, 1.667544729E9, 1.667544777E9, 1.667544825E9, 1.667544873E9, 1.667544921E9, 1.667544969E9, 1.667545017E9, 1.667545065E9, 1.667545113E9, 1.667545161E9, 1.667545209E9, 1.667545257E9, 1.667545305E9, 1.667545353E9, 1.667545401E9, 1.667545449E9, 1.667545497E9, 1.667545545E9, 1.667545593E9, 1.667545641E9, 1.667545689E9, 1.667545737E9, 1.667545785E9, 1.667545833E9, 1.667545881E9, 1.667545929E9, 1.667545977E9, 1.667546025E9, 1.667546073E9, 1.667546121E9, 1.667546169E9, 1.667546217E9, 1.667546265E9, 1.667546313E9, 1.667546361E9, 1.667546409E9, 1.667546457E9, 1.667546505E9, 1.667546553E9, 1.667546601E9, 1.667546649E9, 1.667546697E9, 1.667546745E9, 1.667546793E9, 1.667546841E9, 1.667546889E9, 1.667546937E9, 1.667546985E9, 1.667547033E9, 1.667547081E9, 1.667547129E9, 1.667547177E9, 1.667547225E9, 1.667547273E9, 1.667547321E9, 1.667547369E9, 1.66754772E9, 1.6675479E9, 1.667553492E9, 1.66755354E9, 1.667553588E9, 1.667553636E9, 1.667553684E9, 1.667553732E9, 1.66755378E9, 1.667553828E9, 1.667553876E9, 1.667553924E9, 1.667553972E9, 1.66755402E9, 1.667554068E9, 1.667554116E9, 1.667554164E9, 1.667554212E9, 1.66755426E9, 1.667554308E9, 1.667554356E9, 1.667554404E9, 1.667554452E9, 1.6675545E9, 1.667554548E9, 1.667554596E9, 1.667554644E9, 1.667554692E9, 1.66755474E9, 1.667554788E9, 1.667554836E9, 1.667554884E9, 1.667554932E9, 1.66755498E9, 1.667555028E9, 1.667555076E9, 1.667555124E9, 1.667555172E9, 1.66755522E9, 1.667555268E9, 1.667555316E9, 1.667555364E9, 1.667555412E9, 1.66755546E9, 1.667555508E9, 1.667555556E9, 1.667555604E9, 1.667555652E9, 1.6675557E9, 1.667555748E9, 1.667555796E9, 1.667555844E9, 1.667555892E9, 1.66755594E9, 1.667555988E9, 1.667556036E9, 1.667556084E9, 1.667556132E9, 1.66755618E9, 1.667556228E9, 1.667556276E9, 1.667556324E9, 1.667556372E9, 1.66755642E9, 1.667556468E9, 1.667556516E9, 1.667556564E9, 1.667556612E9, 1.66755666E9, 1.667556708E9, 1.667556756E9, 1.667556804E9, 1.667556852E9, 1.6675569E9, 1.66755726E9, 1.66755744E9, 1.667563171E9, 1.667563219E9, 1.667563267E9, 1.667563315E9, 1.667563363E9, 1.667563411E9, 1.667563459E9, 1.667563507E9, 1.667563555E9, 1.667563603E9, 1.667563651E9, 1.667563699E9, 1.667563747E9, 1.667563795E9, 1.667563843E9, 1.667563891E9, 1.667563939E9, 1.667563987E9, 1.667564035E9, 1.667564083E9, 1.667564131E9, 1.667564179E9, 1.667564227E9, 1.667564275E9, 1.667564323E9, 1.667564371E9, 1.667564419E9, 1.667564467E9, 1.667564515E9, 1.667564563E9, 1.667564611E9, 1.667564659E9, 1.667564707E9, 1.667564755E9, 1.667564803E9, 1.667564851E9, 1.667564899E9, 1.667564947E9, 1.667564995E9, 1.667565043E9, 1.667565091E9, 1.667565139E9, 1.667565187E9, 1.667565235E9, 1.667565283E9, 1.667565331E9, 1.667565379E9, 1.667565427E9, 1.667565475E9, 1.667565523E9, 1.667565571E9, 1.667565619E9, 1.667565667E9, 1.667565715E9, 1.667565763E9, 1.667565811E9, 1.667565859E9, 1.667565907E9, 1.667565955E9, 1.667566003E9, 1.667566051E9, 1.667566099E9, 1.667566147E9, 1.667566195E9, 1.667566243E9, 1.667566291E9, 1.667566339E9, 1.66756662E9, 1.6675668E9, 1.667572468E9, 1.667572516E9, 1.667572564E9, 1.667572612E9, 1.66757266E9, 1.667572708E9, 1.667572756E9, 1.667572804E9, 1.667572852E9, 1.6675729E9, 1.667572948E9, 1.667572996E9, 1.667573044E9, 1.667573092E9, 1.66757314E9, 1.667573188E9, 1.667573236E9, 1.667573284E9, 1.667573332E9, 1.66757338E9, 1.667573428E9, 1.667573476E9, 1.667573524E9, 1.667573572E9, 1.66757362E9, 1.667573668E9, 1.667573716E9, 1.667573764E9, 1.667573812E9, 1.66757386E9, 1.667573908E9, 1.667573956E9, 1.667574004E9, 1.667574052E9, 1.6675741E9, 1.667574148E9, 1.667574196E9, 1.667574244E9, 1.667574292E9, 1.66757434E9, 1.667574388E9, 1.667574436E9, 1.667574484E9, 1.667574532E9, 1.66757458E9, 1.667574628E9, 1.667574676E9, 1.667574724E9, 1.667574772E9, 1.66757482E9, 1.667574868E9, 1.667574916E9, 1.667574964E9, 1.667575012E9, 1.66757506E9, 1.667575108E9, 1.667575156E9, 1.667575204E9, 1.667575252E9, 1.6675753E9, 1.667575348E9, 1.667575396E9, 1.667575444E9, 1.667575492E9, 1.66757554E9, 1.667575588E9, 1.667575636E9, 1.667575684E9, 1.667575732E9, 1.66757578E9, 1.66757616E9, 1.66757634E9, 1.667581918E9, 1.667581966E9, 1.667582014E9, 1.667582062E9, 1.66758211E9, 1.667582158E9, 1.667582206E9, 1.667582254E9, 1.667582302E9, 1.66758235E9, 1.667582398E9, 1.667582446E9, 1.667582494E9, 1.667582542E9, 1.66758259E9, 1.667582638E9, 1.667582686E9, 1.667582734E9, 1.667582782E9, 1.66758283E9, 1.667582878E9, 1.667582926E9, 1.667582974E9, 1.667583022E9, 1.66758307E9, 1.667583118E9, 1.667583166E9, 1.667583214E9, 1.667583262E9, 1.66758331E9, 1.667583358E9, 1.667583406E9, 1.667583454E9, 1.667583502E9, 1.66758355E9, 1.667583598E9, 1.667583646E9, 1.667583694E9, 1.667583742E9, 1.66758379E9, 1.667583838E9, 1.667583886E9, 1.667583934E9, 1.667583982E9, 1.66758403E9, 1.667584078E9, 1.667584126E9, 1.667584174E9, 1.667584222E9, 1.66758427E9, 1.667584318E9, 1.667584366E9, 1.667584414E9, 1.667584462E9, 1.66758451E9, 1.667584558E9, 1.667584606E9, 1.667584654E9, 1.667584702E9, 1.66758475E9, 1.667584798E9, 1.667584846E9, 1.667584894E9, 1.667584942E9, 1.66758499E9, 1.667585038E9, 1.667585086E9, 1.667585134E9, 1.667585182E9, 1.66758523E9, 1.66758558E9, 1.66758576E9, 1.667591371E9, 1.667591419E9, 1.667591467E9, 1.667591515E9, 1.667591563E9, 1.667591611E9, 1.667591659E9, 1.667591707E9, 1.667591755E9, 1.667591803E9, 1.667591851E9, 1.667591899E9, 1.667591947E9, 1.667591995E9, 1.667592043E9, 1.667592091E9, 1.667592139E9, 1.667592187E9, 1.667592235E9, 1.667592283E9, 1.667592331E9, 1.667592379E9, 1.667592427E9, 1.667592475E9, 1.667592523E9, 1.667592571E9, 1.667592619E9, 1.667592667E9, 1.667592715E9, 1.667592763E9, 1.667592811E9, 1.667592859E9, 1.667592907E9, 1.667592955E9, 1.667593003E9, 1.667593051E9, 1.667593099E9, 1.667593147E9, 1.667593195E9, 1.667593243E9, 1.667593291E9, 1.667593339E9, 1.667593387E9, 1.667593435E9, 1.667593483E9, 1.667593531E9, 1.667593579E9, 1.667593627E9, 1.667593675E9, 1.667593723E9, 1.667593771E9, 1.667593819E9, 1.667593867E9, 1.667593915E9, 1.667593963E9, 1.667594011E9, 1.667594059E9, 1.667594107E9, 1.667594155E9, 1.667594203E9, 1.667594251E9, 1.667594299E9, 1.667594347E9, 1.667594395E9, 1.667594443E9, 1.667594491E9, 1.667594539E9, 1.66759482E9, 1.66759494E9, 1.66760064E9, 1.667600688E9, 1.667600736E9, 1.667600784E9, 1.667600832E9, 1.66760088E9, 1.667600928E9, 1.667600976E9, 1.667601024E9, 1.667601072E9, 1.66760112E9, 1.667601168E9, 1.667601216E9, 1.667601264E9, 1.667601312E9, 1.66760136E9, 1.667601408E9, 1.667601456E9, 1.667601504E9, 1.667601552E9, 1.6676016E9, 1.667601648E9, 1.667601696E9, 1.667601744E9, 1.667601792E9, 1.66760184E9, 1.667601888E9, 1.667601936E9, 1.667601984E9, 1.667602032E9, 1.66760208E9, 1.667602128E9, 1.667602176E9, 1.667602224E9, 1.667602272E9, 1.66760232E9, 1.667602368E9, 1.667602416E9, 1.667602464E9, 1.667602512E9, 1.66760256E9, 1.667602608E9, 1.667602656E9, 1.667602704E9, 1.667602752E9, 1.6676028E9, 1.667602848E9, 1.667602896E9, 1.667602944E9, 1.667602992E9, 1.66760304E9, 1.667603088E9, 1.667603136E9, 1.667603184E9, 1.667603232E9, 1.66760328E9, 1.667603328E9, 1.667603376E9, 1.667603424E9, 1.667603472E9, 1.66760352E9, 1.667603568E9, 1.667603616E9, 1.667603664E9, 1.667603712E9, 1.66760376E9, 1.667603808E9, 1.667603856E9, 1.667603904E9, 1.667603952E9, 1.667604E9, 1.6676043E9, 1.66760448E9, 1.667610334E9, 1.667610382E9, 1.66761043E9, 1.667610478E9, 1.667610526E9, 1.667610574E9, 1.667610622E9, 1.66761067E9, 1.667610718E9, 1.667610766E9, 1.667610814E9, 1.667610862E9, 1.66761091E9, 1.667610958E9, 1.667611006E9, 1.667611054E9, 1.667611102E9, 1.66761115E9, 1.667611198E9, 1.667611246E9, 1.667611294E9, 1.667611342E9, 1.66761139E9, 1.667611438E9, 1.667611486E9, 1.667611534E9, 1.667611582E9, 1.66761163E9, 1.667611678E9, 1.667611726E9, 1.667611774E9, 1.667611822E9, 1.66761187E9, 1.667611918E9, 1.667611966E9, 1.667612014E9, 1.667612062E9, 1.66761211E9, 1.667612158E9, 1.667612206E9, 1.667612254E9, 1.667612302E9, 1.66761235E9, 1.667612398E9, 1.667612446E9, 1.667612494E9, 1.667612542E9, 1.66761259E9, 1.667612638E9, 1.667612686E9, 1.667612734E9, 1.667612782E9, 1.66761283E9, 1.667612878E9, 1.667612926E9, 1.667612974E9, 1.667613022E9, 1.66761307E9, 1.667613118E9, 1.667613166E9, 1.667613214E9, 1.667613262E9, 1.66761331E9, 1.667613358E9, 1.667613406E9, 1.667613454E9, 1.667613502E9, 1.66761355E9, 1.667613598E9, 1.667613646E9, 1.667613694E9, 1.667613742E9, 1.66761379E9, 1.66761414E9, 1.66761432E9, 1.667620017E9, 1.667620065E9, 1.667620113E9, 1.667620161E9, 1.667620209E9, 1.667620257E9, 1.667620305E9, 1.667620353E9, 1.667620401E9, 1.667620449E9, 1.667620497E9, 1.667620545E9, 1.667620593E9, 1.667620641E9, 1.667620689E9, 1.667620737E9, 1.667620785E9, 1.667620833E9, 1.667620881E9, 1.667620929E9, 1.667620977E9, 1.667621025E9, 1.667621073E9, 1.667621121E9, 1.667621169E9, 1.667621217E9, 1.667621265E9, 1.667621313E9, 1.667621361E9, 1.667621409E9, 1.667621457E9, 1.667621505E9, 1.667621553E9, 1.667621601E9, 1.667621649E9, 1.667621697E9, 1.667621745E9, 1.667621793E9, 1.667621841E9, 1.667621889E9, 1.667621937E9, 1.667621985E9, 1.667622033E9, 1.667622081E9, 1.667622129E9, 1.667622177E9, 1.667622225E9, 1.667622273E9, 1.667622321E9, 1.667622369E9, 1.667622417E9, 1.667622465E9, 1.667622513E9, 1.667622561E9, 1.667622609E9, 1.667622657E9, 1.667622705E9, 1.667622753E9, 1.667622801E9, 1.667622849E9, 1.667622897E9, 1.667622945E9, 1.667622993E9, 1.667623041E9, 1.667623089E9, 1.667623137E9, 1.667623185E9, 1.667623233E9, 1.667623281E9, 1.667623329E9, 1.66762362E9, 1.6676238E9, 1.667629451E9, 1.667629499E9, 1.667629547E9, 1.667629595E9, 1.667629643E9, 1.667629691E9, 1.667629739E9, 1.667629787E9, 1.667629835E9, 1.667629883E9, 1.667629931E9, 1.667629979E9, 1.667630027E9, 1.667630075E9, 1.667630123E9, 1.667630171E9, 1.667630219E9, 1.667630267E9, 1.667630315E9, 1.667630363E9, 1.667630411E9, 1.667630459E9, 1.667630507E9, 1.667630555E9, 1.667630603E9, 1.667630651E9, 1.667630699E9, 1.667630747E9, 1.667630795E9, 1.667630843E9, 1.667630891E9, 1.667630939E9, 1.667630987E9, 1.667631035E9, 1.667631083E9, 1.667631131E9, 1.667631179E9, 1.667631227E9, 1.667631275E9, 1.667631323E9, 1.667631371E9, 1.667631419E9, 1.667631467E9, 1.667631515E9, 1.667631563E9, 1.667631611E9, 1.667631659E9, 1.667631707E9, 1.667631755E9, 1.667631803E9, 1.667631851E9, 1.667631899E9, 1.667631947E9, 1.667631995E9, 1.667632043E9, 1.667632091E9, 1.667632139E9, 1.667632187E9, 1.667632235E9, 1.667632283E9, 1.667632331E9, 1.667632379E9, 1.667632427E9, 1.667632475E9, 1.667632523E9, 1.667632571E9, 1.667632619E9, 1.66763292E9, 1.6676331E9, 1.667638814E9, 1.667638862E9, 1.66763891E9, 1.667638958E9, 1.667639006E9, 1.667639054E9, 1.667639102E9, 1.66763915E9, 1.667639198E9, 1.667639246E9, 1.667639294E9, 1.667639342E9, 1.66763939E9, 1.667639438E9, 1.667639486E9, 1.667639534E9, 1.667639582E9, 1.66763963E9, 1.667639678E9, 1.667639726E9, 1.667639774E9, 1.667639822E9, 1.66763987E9, 1.667639918E9, 1.667639966E9, 1.667640014E9, 1.667640062E9, 1.66764011E9, 1.667640158E9, 1.667640206E9, 1.667640254E9, 1.667640302E9, 1.66764035E9, 1.667640398E9, 1.667640446E9, 1.667640494E9, 1.667640542E9, 1.66764059E9, 1.667640638E9, 1.667640686E9, 1.667640734E9, 1.667640782E9, 1.66764083E9, 1.667640878E9, 1.667640926E9, 1.667640974E9, 1.667641022E9, 1.66764107E9, 1.667641118E9, 1.667641166E9, 1.667641214E9, 1.667641262E9, 1.66764131E9, 1.667641358E9, 1.667641406E9, 1.667641454E9, 1.667641502E9, 1.66764155E9, 1.667641598E9, 1.667641646E9, 1.667641694E9, 1.667641742E9, 1.66764179E9, 1.667641838E9, 1.667641886E9, 1.667641934E9, 1.667641982E9, 1.66764203E9, 1.66764234E9, 1.66764252E9, 1.667648246E9, 1.667648294E9, 1.667648342E9, 1.66764839E9, 1.667648438E9, 1.667648486E9, 1.667648534E9, 1.667648582E9, 1.66764863E9, 1.667648678E9, 1.667648726E9, 1.667648774E9, 1.667648822E9, 1.66764887E9, 1.667648918E9, 1.667648966E9, 1.667649014E9, 1.667649062E9, 1.66764911E9, 1.667649158E9, 1.667649206E9, 1.667649254E9, 1.667649302E9, 1.66764935E9, 1.667649398E9, 1.667649446E9, 1.667649494E9, 1.667649542E9, 1.66764959E9, 1.667649638E9, 1.667649686E9, 1.667649734E9, 1.667649782E9, 1.66764983E9, 1.667649878E9, 1.667649926E9, 1.667649974E9, 1.667650022E9, 1.66765007E9, 1.667650118E9, 1.667650166E9, 1.667650214E9, 1.667650262E9, 1.66765031E9, 1.667650358E9, 1.667650406E9, 1.667650454E9, 1.667650502E9, 1.66765055E9, 1.667650598E9, 1.667650646E9, 1.667650694E9, 1.667650742E9, 1.66765079E9, 1.667650838E9, 1.667650886E9, 1.667650934E9, 1.667650982E9, 1.66765103E9, 1.667651078E9, 1.667651126E9, 1.667651174E9, 1.667651222E9, 1.66765127E9, 1.667651318E9, 1.667651366E9, 1.667651414E9, 1.667651462E9, 1.66765151E9, 1.66765188E9, 1.667652E9, 1.667657672E9, 1.66765772E9, 1.667657768E9, 1.667657816E9, 1.667657864E9, 1.667657912E9, 1.66765796E9, 1.667658008E9, 1.667658056E9, 1.667658104E9, 1.667658152E9, 1.6676582E9, 1.667658248E9, 1.667658296E9, 1.667658344E9, 1.667658392E9, 1.66765844E9, 1.667658488E9, 1.667658536E9, 1.667658584E9, 1.667658632E9, 1.66765868E9, 1.667658728E9, 1.667658776E9, 1.667658824E9, 1.667658872E9, 1.66765892E9, 1.667658968E9, 1.667659016E9, 1.667659064E9, 1.667659112E9, 1.66765916E9, 1.667659208E9, 1.667659256E9, 1.667659304E9, 1.667659352E9, 1.6676594E9, 1.667659448E9, 1.667659496E9, 1.667659544E9, 1.667659592E9, 1.66765964E9, 1.667659688E9, 1.667659736E9, 1.667659784E9, 1.667659832E9, 1.66765988E9, 1.667659928E9, 1.667659976E9, 1.667660024E9, 1.667660072E9, 1.66766012E9, 1.667660168E9, 1.667660216E9, 1.667660264E9, 1.667660312E9, 1.66766036E9, 1.667660408E9, 1.667660456E9, 1.667660504E9, 1.667660552E9, 1.6676606E9, 1.667660648E9, 1.667660696E9, 1.667660744E9, 1.667660792E9, 1.66766084E9, 1.667660888E9, 1.667660936E9, 1.667660984E9, 1.667661032E9, 1.66766108E9, 1.66766136E9, 1.66766154E9, 1.667667297E9, 1.667667345E9, 1.667667393E9, 1.667667441E9, 1.667667489E9, 1.667667537E9, 1.667667585E9, 1.667667633E9, 1.667667681E9, 1.667667729E9, 1.667667777E9, 1.667667825E9, 1.667667873E9, 1.667667921E9, 1.667667969E9, 1.667668017E9, 1.667668065E9, 1.667668113E9, 1.667668161E9, 1.667668209E9, 1.667668257E9, 1.667668305E9, 1.667668353E9, 1.667668401E9, 1.667668449E9, 1.667668497E9, 1.667668545E9, 1.667668593E9, 1.667668641E9, 1.667668689E9, 1.667668737E9, 1.667668785E9, 1.667668833E9, 1.667668881E9, 1.667668929E9, 1.667668977E9, 1.667669025E9, 1.667669073E9, 1.667669121E9, 1.667669169E9, 1.667669217E9, 1.667669265E9, 1.667669313E9, 1.667669361E9, 1.667669409E9, 1.667669457E9, 1.667669505E9, 1.667669553E9, 1.667669601E9, 1.667669649E9, 1.667669697E9, 1.667669745E9, 1.667669793E9, 1.667669841E9, 1.667669889E9, 1.667669937E9, 1.667669985E9, 1.667670033E9, 1.667670081E9, 1.667670129E9, 1.667670177E9, 1.667670225E9, 1.667670273E9, 1.667670321E9, 1.667670369E9, 1.667670417E9, 1.667670465E9, 1.667670513E9, 1.667670561E9, 1.667670609E9, 1.6676709E9, 1.66767108E9, 1.667676687E9, 1.667676735E9, 1.667676783E9, 1.667676831E9, 1.667676879E9, 1.667676927E9, 1.667676975E9, 1.667677023E9, 1.667677071E9, 1.667677119E9, 1.667677167E9, 1.667677215E9, 1.667677263E9, 1.667677311E9, 1.667677359E9, 1.667677407E9, 1.667677455E9, 1.667677503E9, 1.667677551E9, 1.667677599E9, 1.667677647E9, 1.667677695E9, 1.667677743E9, 1.667677791E9, 1.667677839E9, 1.667677887E9, 1.667677935E9, 1.667677983E9, 1.667678031E9, 1.667678079E9, 1.667678127E9, 1.667678175E9, 1.667678223E9, 1.667678271E9, 1.667678319E9, 1.667678367E9, 1.667678415E9, 1.667678463E9, 1.667678511E9, 1.667678559E9, 1.667678607E9, 1.667678655E9, 1.667678703E9, 1.667678751E9, 1.667678799E9, 1.667678847E9, 1.667678895E9, 1.667678943E9, 1.667678991E9, 1.667679039E9, 1.667679087E9, 1.667679135E9, 1.667679183E9, 1.667679231E9, 1.667679279E9, 1.667679327E9, 1.667679375E9, 1.667679423E9, 1.667679471E9, 1.667679519E9, 1.667679567E9, 1.667679615E9, 1.667679663E9, 1.667679711E9, 1.667679759E9, 1.667679807E9, 1.667679855E9, 1.667679903E9, 1.667679951E9, 1.667679999E9, 1.66768038E9, 1.66768056E9, 1.667686333E9, 1.667686381E9, 1.667686429E9, 1.667686477E9, 1.667686525E9, 1.667686573E9, 1.667686621E9, 1.667686669E9, 1.667686717E9, 1.667686765E9, 1.667686813E9, 1.667686861E9, 1.667686909E9, 1.667686957E9, 1.667687005E9, 1.667687053E9, 1.667687101E9, 1.667687149E9, 1.667687197E9, 1.667687245E9, 1.667687293E9, 1.667687341E9, 1.667687389E9, 1.667687437E9, 1.667687485E9, 1.667687533E9, 1.667687581E9, 1.667687629E9, 1.667687677E9, 1.667687725E9, 1.667687773E9, 1.667687821E9, 1.667687869E9, 1.667687917E9, 1.667687965E9, 1.667688013E9, 1.667688061E9, 1.667688109E9, 1.667688157E9, 1.667688205E9, 1.667688253E9, 1.667688301E9, 1.667688349E9, 1.667688397E9, 1.667688445E9, 1.667688493E9, 1.667688541E9, 1.667688589E9, 1.667688637E9, 1.667688685E9, 1.667688733E9, 1.667688781E9, 1.667688829E9, 1.667688877E9, 1.667688925E9, 1.667688973E9, 1.667689021E9, 1.667689069E9, 1.667689117E9, 1.667689165E9, 1.667689213E9, 1.667689261E9, 1.667689309E9, 1.667689357E9, 1.667689405E9, 1.667689453E9, 1.667689501E9, 1.667689549E9, 1.6676898E9, 1.66768998E9, 1.667695669E9, 1.667695717E9, 1.667695765E9, 1.667695813E9, 1.667695861E9, 1.667695909E9, 1.667695957E9, 1.667696005E9, 1.667696053E9, 1.667696101E9, 1.667696149E9, 1.667696197E9, 1.667696245E9, 1.667696293E9, 1.667696341E9, 1.667696389E9, 1.667696437E9, 1.667696485E9, 1.667696533E9, 1.667696581E9, 1.667696629E9, 1.667696677E9, 1.667696725E9, 1.667696773E9, 1.667696821E9, 1.667696869E9, 1.667696917E9, 1.667696965E9, 1.667697013E9, 1.667697061E9, 1.667697109E9, 1.667697157E9, 1.667697205E9, 1.667697253E9, 1.667697301E9, 1.667697349E9, 1.667697397E9, 1.667697445E9, 1.667697493E9, 1.667697541E9, 1.667697589E9, 1.667697637E9, 1.667697685E9, 1.667697733E9, 1.667697781E9, 1.667697829E9, 1.667697877E9, 1.667697925E9, 1.667697973E9, 1.667698021E9, 1.667698069E9, 1.667698117E9, 1.667698165E9, 1.667698213E9, 1.667698261E9, 1.667698309E9, 1.667698357E9, 1.667698405E9, 1.667698453E9, 1.667698501E9, 1.667698549E9, 1.667698597E9, 1.667698645E9, 1.667698693E9, 1.667698741E9, 1.667698789E9, 1.667698837E9, 1.667698885E9, 1.667698933E9, 1.667698981E9, 1.667699029E9, 1.6676994E9, 1.66769964E9, 1.66770524E9, 1.667705288E9, 1.667705336E9, 1.667705384E9, 1.667705432E9, 1.66770548E9, 1.667705528E9, 1.667705576E9, 1.667705624E9, 1.667705672E9, 1.66770572E9, 1.667705768E9, 1.667705816E9, 1.667705864E9, 1.667705912E9, 1.66770596E9, 1.667706008E9, 1.667706056E9, 1.667706104E9, 1.667706152E9, 1.6677062E9, 1.667706248E9, 1.667706296E9, 1.667706344E9, 1.667706392E9, 1.66770644E9, 1.667706488E9, 1.667706536E9, 1.667706584E9, 1.667706632E9, 1.66770668E9, 1.667706728E9, 1.667706776E9, 1.667706824E9, 1.667706872E9, 1.66770692E9, 1.667706968E9, 1.667707016E9, 1.667707064E9, 1.667707112E9, 1.66770716E9, 1.667707208E9, 1.667707256E9, 1.667707304E9, 1.667707352E9, 1.6677074E9, 1.667707448E9, 1.667707496E9, 1.667707544E9, 1.667707592E9, 1.66770764E9, 1.667707688E9, 1.667707736E9, 1.667707784E9, 1.667707832E9, 1.66770788E9, 1.667707928E9, 1.667707976E9, 1.667708024E9, 1.667708072E9, 1.66770812E9, 1.667708168E9, 1.667708216E9, 1.667708264E9, 1.667708312E9, 1.66770836E9, 1.667708408E9, 1.667708456E9, 1.667708504E9, 1.667708552E9, 1.6677086E9, 1.66770894E9, 1.66770912E9, 1.667714834E9, 1.667714882E9, 1.66771493E9, 1.667714978E9, 1.667715026E9, 1.667715074E9, 1.667715122E9, 1.66771517E9, 1.667715218E9, 1.667715266E9, 1.667715314E9, 1.667715362E9, 1.66771541E9, 1.667715458E9, 1.667715506E9, 1.667715554E9, 1.667715602E9, 1.66771565E9, 1.667715698E9, 1.667715746E9, 1.667715794E9, 1.667715842E9, 1.66771589E9, 1.667715938E9, 1.667715986E9, 1.667716034E9, 1.667716082E9, 1.66771613E9, 1.667716178E9, 1.667716226E9, 1.667716274E9, 1.667716322E9, 1.66771637E9, 1.667716418E9, 1.667716466E9, 1.667716514E9, 1.667716562E9, 1.66771661E9, 1.667716658E9, 1.667716706E9, 1.667716754E9, 1.667716802E9, 1.66771685E9, 1.667716898E9, 1.667716946E9, 1.667716994E9, 1.667717042E9, 1.66771709E9, 1.667717138E9, 1.667717186E9, 1.667717234E9, 1.667717282E9, 1.66771733E9, 1.667717378E9, 1.667717426E9, 1.667717474E9, 1.667717522E9, 1.66771757E9, 1.667717618E9, 1.667717666E9, 1.667717714E9, 1.667717762E9, 1.66771781E9, 1.667717858E9, 1.667717906E9, 1.667717954E9, 1.667718002E9, 1.66771805E9, 1.66771842E9, 1.6677186E9, 1.66772424E9, 1.667724288E9, 1.667724336E9, 1.667724384E9, 1.667724432E9, 1.66772448E9, 1.667724528E9, 1.667724576E9, 1.667724624E9, 1.667724672E9, 1.66772472E9, 1.667724768E9, 1.667724816E9, 1.667724864E9, 1.667724912E9, 1.66772496E9, 1.667725008E9, 1.667725056E9, 1.667725104E9, 1.667725152E9, 1.6677252E9, 1.667725248E9, 1.667725296E9, 1.667725344E9, 1.667725392E9, 1.66772544E9, 1.667725488E9, 1.667725536E9, 1.667725584E9, 1.667725632E9, 1.66772568E9, 1.667725728E9, 1.667725776E9, 1.667725824E9, 1.667725872E9, 1.66772592E9, 1.667725968E9, 1.667726016E9, 1.667726064E9, 1.667726112E9, 1.66772616E9, 1.667726208E9, 1.667726256E9, 1.667726304E9, 1.667726352E9, 1.6677264E9, 1.667726448E9, 1.667726496E9, 1.667726544E9, 1.667726592E9, 1.66772664E9, 1.667726688E9, 1.667726736E9, 1.667726784E9, 1.667726832E9, 1.66772688E9, 1.667726928E9, 1.667726976E9, 1.667727024E9, 1.667727072E9, 1.66772712E9, 1.667727168E9, 1.667727216E9, 1.667727264E9, 1.667727312E9, 1.66772736E9, 1.667727408E9, 1.667727456E9, 1.667727504E9, 1.667727552E9, 1.6677276E9, 1.6677279E9, 1.66772808E9, 1.667733646E9, 1.667733694E9, 1.667733742E9, 1.66773379E9, 1.667733838E9, 1.667733886E9, 1.667733934E9, 1.667733982E9, 1.66773403E9, 1.667734078E9, 1.667734126E9, 1.667734174E9, 1.667734222E9, 1.66773427E9, 1.667734318E9, 1.667734366E9, 1.667734414E9, 1.667734462E9, 1.66773451E9, 1.667734558E9, 1.667734606E9, 1.667734654E9, 1.667734702E9, 1.66773475E9, 1.667734798E9, 1.667734846E9, 1.667734894E9, 1.667734942E9, 1.66773499E9, 1.667735038E9, 1.667735086E9, 1.667735134E9, 1.667735182E9, 1.66773523E9, 1.667735278E9, 1.667735326E9, 1.667735374E9, 1.667735422E9, 1.66773547E9, 1.667735518E9, 1.667735566E9, 1.667735614E9, 1.667735662E9, 1.66773571E9, 1.667735758E9, 1.667735806E9, 1.667735854E9, 1.667735902E9, 1.66773595E9, 1.667735998E9, 1.667736046E9, 1.667736094E9, 1.667736142E9, 1.66773619E9, 1.667736238E9, 1.667736286E9, 1.667736334E9, 1.667736382E9, 1.66773643E9, 1.667736478E9, 1.667736526E9, 1.667736574E9, 1.667736622E9, 1.66773667E9, 1.667736718E9, 1.667736766E9, 1.667736814E9, 1.667736862E9, 1.66773691E9, 1.66773732E9, 1.66773744E9, 1.667743087E9, 1.667743135E9, 1.667743183E9, 1.667743231E9, 1.667743279E9, 1.667743327E9, 1.667743375E9, 1.667743423E9, 1.667743471E9, 1.667743519E9, 1.667743567E9, 1.667743615E9, 1.667743663E9, 1.667743711E9, 1.667743759E9, 1.667743807E9, 1.667743855E9, 1.667743903E9, 1.667743951E9, 1.667743999E9, 1.667744047E9, 1.667744095E9, 1.667744143E9, 1.667744191E9, 1.667744239E9, 1.667744287E9, 1.667744335E9, 1.667744383E9, 1.667744431E9, 1.667744479E9, 1.667744527E9, 1.667744575E9, 1.667744623E9, 1.667744671E9, 1.667744719E9, 1.667744767E9, 1.667744815E9, 1.667744863E9, 1.667744911E9, 1.667744959E9, 1.667745007E9, 1.667745055E9, 1.667745103E9, 1.667745151E9, 1.667745199E9, 1.667745247E9, 1.667745295E9, 1.667745343E9, 1.667745391E9, 1.667745439E9, 1.667745487E9, 1.667745535E9, 1.667745583E9, 1.667745631E9, 1.667745679E9, 1.667745727E9, 1.667745775E9, 1.667745823E9, 1.667745871E9, 1.667745919E9, 1.667745967E9, 1.667746015E9, 1.667746063E9, 1.667746111E9, 1.667746159E9, 1.667746207E9, 1.667746255E9, 1.667746303E9, 1.667746351E9, 1.667746399E9, 1.66774668E9, 1.66774686E9, 1.667752465E9, 1.667752513E9, 1.667752561E9, 1.667752609E9, 1.667752657E9, 1.667752705E9, 1.667752753E9, 1.667752801E9, 1.667752849E9, 1.667752897E9, 1.667752945E9, 1.667752993E9, 1.667753041E9, 1.667753089E9, 1.667753137E9, 1.667753185E9, 1.667753233E9, 1.667753281E9, 1.667753329E9, 1.667753377E9, 1.667753425E9, 1.667753473E9, 1.667753521E9, 1.667753569E9, 1.667753617E9, 1.667753665E9, 1.667753713E9, 1.667753761E9, 1.667753809E9, 1.667753857E9, 1.667753905E9, 1.667753953E9, 1.667754001E9, 1.667754049E9, 1.667754097E9, 1.667754145E9, 1.667754193E9, 1.667754241E9, 1.667754289E9, 1.667754337E9, 1.667754385E9, 1.667754433E9, 1.667754481E9, 1.667754529E9, 1.667754577E9, 1.667754625E9, 1.667754673E9, 1.667754721E9, 1.667754769E9, 1.667754817E9, 1.667754865E9, 1.667754913E9, 1.667754961E9, 1.667755009E9, 1.667755057E9, 1.667755105E9, 1.667755153E9, 1.667755201E9, 1.667755249E9, 1.667755297E9, 1.667755345E9, 1.667755393E9, 1.667755441E9, 1.667755489E9, 1.667755537E9, 1.667755585E9, 1.667755633E9, 1.667755681E9, 1.667755729E9, 1.66775598E9, 1.66775616E9, 1.667761744E9, 1.667761792E9, 1.66776184E9, 1.667761888E9, 1.667761936E9, 1.667761984E9, 1.667762032E9, 1.66776208E9, 1.667762128E9, 1.667762176E9, 1.667762224E9, 1.667762272E9, 1.66776232E9, 1.667762368E9, 1.667762416E9, 1.667762464E9, 1.667762512E9, 1.66776256E9, 1.667762608E9, 1.667762656E9, 1.667762704E9, 1.667762752E9, 1.6677628E9, 1.667762848E9, 1.667762896E9, 1.667762944E9, 1.667762992E9, 1.66776304E9, 1.667763088E9, 1.667763136E9, 1.667763184E9, 1.667763232E9, 1.66776328E9, 1.667763328E9, 1.667763376E9, 1.667763424E9, 1.667763472E9, 1.66776352E9, 1.667763568E9, 1.667763616E9, 1.667763664E9, 1.667763712E9, 1.66776376E9, 1.667763808E9, 1.667763856E9, 1.667763904E9, 1.667763952E9, 1.667764E9, 1.667764048E9, 1.667764096E9, 1.667764144E9, 1.667764192E9, 1.66776424E9, 1.667764288E9, 1.667764336E9, 1.667764384E9, 1.667764432E9, 1.66776448E9, 1.667764528E9, 1.667764576E9, 1.667764624E9, 1.667764672E9, 1.66776472E9, 1.667764768E9, 1.667764816E9, 1.667764864E9, 1.667764912E9, 1.66776496E9, 1.66776528E9, 1.66776546E9, 1.667771201E9, 1.667771249E9, 1.667771297E9, 1.667771345E9, 1.667771393E9, 1.667771441E9, 1.667771489E9, 1.667771537E9, 1.667771585E9, 1.667771633E9, 1.667771681E9, 1.667771729E9, 1.667771777E9, 1.667771825E9, 1.667771873E9, 1.667771921E9, 1.667771969E9, 1.667772017E9, 1.667772065E9, 1.667772113E9, 1.667772161E9, 1.667772209E9, 1.667772257E9, 1.667772305E9, 1.667772353E9, 1.667772401E9, 1.667772449E9, 1.667772497E9, 1.667772545E9, 1.667772593E9, 1.667772641E9, 1.667772689E9, 1.667772737E9, 1.667772785E9, 1.667772833E9, 1.667772881E9, 1.667772929E9, 1.667772977E9, 1.667773025E9, 1.667773073E9, 1.667773121E9, 1.667773169E9, 1.667773217E9, 1.667773265E9, 1.667773313E9, 1.667773361E9, 1.667773409E9, 1.667773457E9, 1.667773505E9, 1.667773553E9, 1.667773601E9, 1.667773649E9, 1.667773697E9, 1.667773745E9, 1.667773793E9, 1.667773841E9, 1.667773889E9, 1.667773937E9, 1.667773985E9, 1.667774033E9, 1.667774081E9, 1.667774129E9, 1.667774177E9, 1.667774225E9, 1.667774273E9, 1.667774321E9, 1.667774369E9, 1.667774417E9, 1.667774465E9, 1.667774513E9, 1.667774561E9, 1.667774609E9, 1.66777488E9, 1.66777506E9, 1.667780918E9, 1.667780966E9, 1.667781014E9, 1.667781062E9, 1.66778111E9, 1.667781158E9, 1.667781206E9, 1.667781254E9, 1.667781302E9, 1.66778135E9, 1.667781398E9, 1.667781446E9, 1.667781494E9, 1.667781542E9, 1.66778159E9, 1.667781638E9, 1.667781686E9, 1.667781734E9, 1.667781782E9, 1.66778183E9, 1.667781878E9, 1.667781926E9, 1.667781974E9, 1.667782022E9, 1.66778207E9, 1.667782118E9, 1.667782166E9, 1.667782214E9, 1.667782262E9, 1.66778231E9, 1.667782358E9, 1.667782406E9, 1.667782454E9, 1.667782502E9, 1.66778255E9, 1.667782598E9, 1.667782646E9, 1.667782694E9, 1.667782742E9, 1.66778279E9, 1.667782838E9, 1.667782886E9, 1.667782934E9, 1.667782982E9, 1.66778303E9, 1.667783078E9, 1.667783126E9, 1.667783174E9, 1.667783222E9, 1.66778327E9, 1.667783318E9, 1.667783366E9, 1.667783414E9, 1.667783462E9, 1.66778351E9, 1.667783558E9, 1.667783606E9, 1.667783654E9, 1.667783702E9, 1.66778375E9, 1.667783798E9, 1.667783846E9, 1.667783894E9, 1.667783942E9, 1.66778399E9, 1.667784038E9, 1.667784086E9, 1.667784134E9, 1.667784182E9, 1.66778423E9, 1.66778454E9, 1.66778472E9, 1.667790453E9, 1.667790501E9, 1.667790549E9, 1.667790597E9, 1.667790645E9, 1.667790693E9, 1.667790741E9, 1.667790789E9, 1.667790837E9, 1.667790885E9, 1.667790933E9, 1.667790981E9, 1.667791029E9, 1.667791077E9, 1.667791125E9, 1.667791173E9, 1.667791221E9, 1.667791269E9, 1.667791317E9, 1.667791365E9, 1.667791413E9, 1.667791461E9, 1.667791509E9, 1.667791557E9, 1.667791605E9, 1.667791653E9, 1.667791701E9, 1.667791749E9, 1.667791797E9, 1.667791845E9, 1.667791893E9, 1.667791941E9, 1.667791989E9, 1.667792037E9, 1.667792085E9, 1.667792133E9, 1.667792181E9, 1.667792229E9, 1.667792277E9, 1.667792325E9, 1.667792373E9, 1.667792421E9, 1.667792469E9, 1.667792517E9, 1.667792565E9, 1.667792613E9, 1.667792661E9, 1.667792709E9, 1.667792757E9, 1.667792805E9, 1.667792853E9, 1.667792901E9, 1.667792949E9, 1.667792997E9, 1.667793045E9, 1.667793093E9, 1.667793141E9, 1.667793189E9, 1.667793237E9, 1.667793285E9, 1.667793333E9, 1.667793381E9, 1.667793429E9, 1.667793477E9, 1.667793525E9, 1.667793573E9, 1.667793621E9, 1.667793669E9, 1.66779396E9, 1.66779414E9, 1.667799761E9, 1.667799809E9, 1.667799857E9, 1.667799905E9, 1.667799953E9, 1.667800001E9, 1.667800049E9, 1.667800097E9, 1.667800145E9, 1.667800193E9, 1.667800241E9, 1.667800289E9, 1.667800337E9, 1.667800385E9, 1.667800433E9, 1.667800481E9, 1.667800529E9, 1.667800577E9, 1.667800625E9, 1.667800673E9, 1.667800721E9, 1.667800769E9, 1.667800817E9, 1.667800865E9, 1.667800913E9, 1.667800961E9, 1.667801009E9, 1.667801057E9, 1.667801105E9, 1.667801153E9, 1.667801201E9, 1.667801249E9, 1.667801297E9, 1.667801345E9, 1.667801393E9, 1.667801441E9, 1.667801489E9, 1.667801537E9, 1.667801585E9, 1.667801633E9, 1.667801681E9, 1.667801729E9, 1.667801777E9, 1.667801825E9, 1.667801873E9, 1.667801921E9, 1.667801969E9, 1.667802017E9, 1.667802065E9, 1.667802113E9, 1.667802161E9, 1.667802209E9, 1.667802257E9, 1.667802305E9, 1.667802353E9, 1.667802401E9, 1.667802449E9, 1.667802497E9, 1.667802545E9, 1.667802593E9, 1.667802641E9, 1.667802689E9, 1.667802737E9, 1.667802785E9, 1.667802833E9, 1.667802881E9, 1.667802929E9, 1.667802977E9, 1.667803025E9, 1.667803073E9, 1.667803121E9, 1.667803169E9, 1.66780356E9, 1.66780374E9, 1.667809395E9, 1.667809443E9, 1.667809491E9, 1.667809539E9, 1.667809587E9, 1.667809635E9, 1.667809683E9, 1.667809731E9, 1.667809779E9, 1.667809827E9, 1.667809875E9, 1.667809923E9, 1.667809971E9, 1.667810019E9, 1.667810067E9, 1.667810115E9, 1.667810163E9, 1.667810211E9, 1.667810259E9, 1.667810307E9, 1.667810355E9, 1.667810403E9, 1.667810451E9, 1.667810499E9, 1.667810547E9, 1.667810595E9, 1.667810643E9, 1.667810691E9, 1.667810739E9, 1.667810787E9, 1.667810835E9, 1.667810883E9, 1.667810931E9, 1.667810979E9, 1.667811027E9, 1.667811075E9, 1.667811123E9, 1.667811171E9, 1.667811219E9, 1.667811267E9, 1.667811315E9, 1.667811363E9, 1.667811411E9, 1.667811459E9, 1.667811507E9, 1.667811555E9, 1.667811603E9, 1.667811651E9, 1.667811699E9, 1.667811747E9, 1.667811795E9, 1.667811843E9, 1.667811891E9, 1.667811939E9, 1.667811987E9, 1.667812035E9, 1.667812083E9, 1.667812131E9, 1.667812179E9, 1.667812227E9, 1.667812275E9, 1.667812323E9, 1.667812371E9, 1.667812419E9, 1.667812467E9, 1.667812515E9, 1.667812563E9, 1.667812611E9, 1.667812659E9, 1.66781298E9, 1.66781316E9, 1.667818935E9, 1.667818983E9, 1.667819031E9, 1.667819079E9, 1.667819127E9, 1.667819175E9, 1.667819223E9, 1.667819271E9, 1.667819319E9, 1.667819367E9, 1.667819415E9, 1.667819463E9, 1.667819511E9, 1.667819559E9, 1.667819607E9, 1.667819655E9, 1.667819703E9, 1.667819751E9, 1.667819799E9, 1.667819847E9, 1.667819895E9, 1.667819943E9, 1.667819991E9, 1.667820039E9, 1.667820087E9, 1.667820135E9, 1.667820183E9, 1.667820231E9, 1.667820279E9, 1.667820327E9, 1.667820375E9, 1.667820423E9, 1.667820471E9, 1.667820519E9, 1.667820567E9, 1.667820615E9, 1.667820663E9, 1.667820711E9, 1.667820759E9, 1.667820807E9, 1.667820855E9, 1.667820903E9, 1.667820951E9, 1.667820999E9, 1.667821047E9, 1.667821095E9, 1.667821143E9, 1.667821191E9, 1.667821239E9, 1.667821287E9, 1.667821335E9, 1.667821383E9, 1.667821431E9, 1.667821479E9, 1.667821527E9, 1.667821575E9, 1.667821623E9, 1.667821671E9, 1.667821719E9, 1.667821767E9, 1.667821815E9, 1.667821863E9, 1.667821911E9, 1.667821959E9, 1.667822007E9, 1.667822055E9, 1.667822103E9, 1.667822151E9, 1.667822199E9, 1.66782258E9, 1.66782276E9, 1.66782853E9, 1.667828578E9, 1.667828626E9, 1.667828674E9, 1.667828722E9, 1.66782877E9, 1.667828818E9, 1.667828866E9, 1.667828914E9, 1.667828962E9, 1.66782901E9, 1.667829058E9, 1.667829106E9, 1.667829154E9, 1.667829202E9, 1.66782925E9, 1.667829298E9, 1.667829346E9, 1.667829394E9, 1.667829442E9, 1.66782949E9, 1.667829538E9, 1.667829586E9, 1.667829634E9, 1.667829682E9, 1.66782973E9, 1.667829778E9, 1.667829826E9, 1.667829874E9, 1.667829922E9, 1.66782997E9, 1.667830018E9, 1.667830066E9, 1.667830114E9, 1.667830162E9, 1.66783021E9, 1.667830258E9, 1.667830306E9, 1.667830354E9, 1.667830402E9, 1.66783045E9, 1.667830498E9, 1.667830546E9, 1.667830594E9, 1.667830642E9, 1.66783069E9, 1.667830738E9, 1.667830786E9, 1.667830834E9, 1.667830882E9, 1.66783093E9, 1.667830978E9, 1.667831026E9, 1.667831074E9, 1.667831122E9, 1.66783117E9, 1.667831218E9, 1.667831266E9, 1.667831314E9, 1.667831362E9, 1.66783141E9, 1.667831458E9, 1.667831506E9, 1.667831554E9, 1.667831602E9, 1.66783165E9, 1.667832E9, 1.66783218E9, 1.667837851E9, 1.667837899E9, 1.667837947E9, 1.667837995E9, 1.667838043E9, 1.667838091E9, 1.667838139E9, 1.667838187E9, 1.667838235E9, 1.667838283E9, 1.667838331E9, 1.667838379E9, 1.667838427E9, 1.667838475E9, 1.667838523E9, 1.667838571E9, 1.667838619E9, 1.667838667E9, 1.667838715E9, 1.667838763E9, 1.667838811E9, 1.667838859E9, 1.667838907E9, 1.667838955E9, 1.667839003E9, 1.667839051E9, 1.667839099E9, 1.667839147E9, 1.667839195E9, 1.667839243E9, 1.667839291E9, 1.667839339E9, 1.667839387E9, 1.667839435E9, 1.667839483E9, 1.667839531E9, 1.667839579E9, 1.667839627E9, 1.667839675E9, 1.667839723E9, 1.667839771E9, 1.667839819E9, 1.667839867E9, 1.667839915E9, 1.667839963E9, 1.667840011E9, 1.667840059E9, 1.667840107E9, 1.667840155E9, 1.667840203E9, 1.667840251E9, 1.667840299E9, 1.667840347E9, 1.667840395E9, 1.667840443E9, 1.667840491E9, 1.667840539E9, 1.667840587E9, 1.667840635E9, 1.667840683E9, 1.667840731E9, 1.667840779E9, 1.667840827E9, 1.667840875E9, 1.667840923E9, 1.667840971E9, 1.667841019E9, 1.667841067E9, 1.667841115E9, 1.667841163E9, 1.667841211E9, 1.667841259E9, 1.66784154E9, 1.66784172E9, 1.667847302E9, 1.66784735E9, 1.667847398E9, 1.667847446E9, 1.667847494E9, 1.667847542E9, 1.66784759E9, 1.667847638E9, 1.667847686E9, 1.667847734E9, 1.667847782E9, 1.66784783E9, 1.667847878E9, 1.667847926E9, 1.667847974E9, 1.667848022E9, 1.66784807E9, 1.667848118E9, 1.667848166E9, 1.667848214E9, 1.667848262E9, 1.66784831E9, 1.667848358E9, 1.667848406E9, 1.667848454E9, 1.667848502E9, 1.66784855E9, 1.667848598E9, 1.667848646E9, 1.667848694E9, 1.667848742E9, 1.66784879E9, 1.667848838E9, 1.667848886E9, 1.667848934E9, 1.667848982E9, 1.66784903E9, 1.667849078E9, 1.667849126E9, 1.667849174E9, 1.667849222E9, 1.66784927E9, 1.667849318E9, 1.667849366E9, 1.667849414E9, 1.667849462E9, 1.66784951E9, 1.667849558E9, 1.667849606E9, 1.667849654E9, 1.667849702E9, 1.66784975E9, 1.667849798E9, 1.667849846E9, 1.667849894E9, 1.667849942E9, 1.66784999E9, 1.667850038E9, 1.667850086E9, 1.667850134E9, 1.667850182E9, 1.66785023E9, 1.667850278E9, 1.667850326E9, 1.667850374E9, 1.667850422E9, 1.66785047E9, 1.66785084E9, 1.66785102E9, 1.667856712E9, 1.66785676E9, 1.667856808E9, 1.667856856E9, 1.667856904E9, 1.667856952E9, 1.667857E9, 1.667857048E9, 1.667857096E9, 1.667857144E9, 1.667857192E9, 1.66785724E9, 1.667857288E9, 1.667857336E9, 1.667857384E9, 1.667857432E9, 1.66785748E9, 1.667857528E9, 1.667857576E9, 1.667857624E9, 1.667857672E9, 1.66785772E9, 1.667857768E9, 1.667857816E9, 1.667857864E9, 1.667857912E9, 1.66785796E9, 1.667858008E9, 1.667858056E9, 1.667858104E9, 1.667858152E9, 1.6678582E9, 1.667858248E9, 1.667858296E9, 1.667858344E9, 1.667858392E9, 1.66785844E9, 1.667858488E9, 1.667858536E9, 1.667858584E9, 1.667858632E9, 1.66785868E9, 1.667858728E9, 1.667858776E9, 1.667858824E9, 1.667858872E9, 1.66785892E9, 1.667858968E9, 1.667859016E9, 1.667859064E9, 1.667859112E9, 1.66785916E9, 1.667859208E9, 1.667859256E9, 1.667859304E9, 1.667859352E9, 1.6678594E9, 1.667859448E9, 1.667859496E9, 1.667859544E9, 1.667859592E9, 1.66785964E9, 1.667859688E9, 1.667859736E9, 1.667859784E9, 1.667859832E9, 1.66785988E9, 1.6678602E9, 1.66786038E9, 1.667866048E9, 1.667866096E9, 1.667866144E9, 1.667866192E9, 1.66786624E9, 1.667866288E9, 1.667866336E9, 1.667866384E9, 1.667866432E9, 1.66786648E9, 1.667866528E9, 1.667866576E9, 1.667866624E9, 1.667866672E9, 1.66786672E9, 1.667866768E9, 1.667866816E9, 1.667866864E9, 1.667866912E9, 1.66786696E9, 1.667867008E9, 1.667867056E9, 1.667867104E9, 1.667867152E9, 1.6678672E9, 1.667867248E9, 1.667867296E9, 1.667867344E9, 1.667867392E9, 1.66786744E9, 1.667867488E9, 1.667867536E9, 1.667867584E9, 1.667867632E9, 1.66786768E9, 1.667867728E9, 1.667867776E9, 1.667867824E9, 1.667867872E9, 1.66786792E9, 1.667867968E9, 1.667868016E9, 1.667868064E9, 1.667868112E9, 1.66786816E9, 1.667868208E9, 1.667868256E9, 1.667868304E9, 1.667868352E9, 1.6678684E9, 1.667868448E9, 1.667868496E9, 1.667868544E9, 1.667868592E9, 1.66786864E9, 1.667868688E9, 1.667868736E9, 1.667868784E9, 1.667868832E9, 1.66786888E9, 1.667868928E9, 1.667868976E9, 1.667869024E9, 1.667869072E9, 1.66786912E9, 1.667869168E9, 1.667869216E9, 1.667869264E9, 1.667869312E9, 1.66786936E9, 1.66786962E9, 1.6678698E9, 1.667875462E9, 1.66787551E9, 1.667875558E9, 1.667875606E9, 1.667875654E9, 1.667875702E9, 1.66787575E9, 1.667875798E9, 1.667875846E9, 1.667875894E9, 1.667875942E9, 1.66787599E9, 1.667876038E9, 1.667876086E9, 1.667876134E9, 1.667876182E9, 1.66787623E9, 1.667876278E9, 1.667876326E9, 1.667876374E9, 1.667876422E9, 1.66787647E9, 1.667876518E9, 1.667876566E9, 1.667876614E9, 1.667876662E9, 1.66787671E9, 1.667876758E9, 1.667876806E9, 1.667876854E9, 1.667876902E9, 1.66787695E9, 1.667876998E9, 1.667877046E9, 1.667877094E9, 1.667877142E9, 1.66787719E9, 1.667877238E9, 1.667877286E9, 1.667877334E9, 1.667877382E9, 1.66787743E9, 1.667877478E9, 1.667877526E9, 1.667877574E9, 1.667877622E9, 1.66787767E9, 1.667877718E9, 1.667877766E9, 1.667877814E9, 1.667877862E9, 1.66787791E9, 1.667877958E9, 1.667878006E9, 1.667878054E9, 1.667878102E9, 1.66787815E9, 1.667878198E9, 1.667878246E9, 1.667878294E9, 1.667878342E9, 1.66787839E9, 1.667878438E9, 1.667878486E9, 1.667878534E9, 1.667878582E9, 1.66787863E9, 1.66787892E9, 1.6678791E9, 1.667885153E9, 1.667885201E9, 1.667885249E9, 1.667885297E9, 1.667885345E9, 1.667885393E9, 1.667885441E9, 1.667885489E9, 1.667885537E9, 1.667885585E9, 1.667885633E9, 1.667885681E9, 1.667885729E9, 1.667885777E9, 1.667885825E9, 1.667885873E9, 1.667885921E9, 1.667885969E9, 1.667886017E9, 1.667886065E9, 1.667886113E9, 1.667886161E9, 1.667886209E9, 1.667886257E9, 1.667886305E9, 1.667886353E9, 1.667886401E9, 1.667886449E9, 1.667886497E9, 1.667886545E9, 1.667886593E9, 1.667886641E9, 1.667886689E9, 1.667886737E9, 1.667886785E9, 1.667886833E9, 1.667886881E9, 1.667886929E9, 1.667886977E9, 1.667887025E9, 1.667887073E9, 1.667887121E9, 1.667887169E9, 1.667887217E9, 1.667887265E9, 1.667887313E9, 1.667887361E9, 1.667887409E9, 1.667887457E9, 1.667887505E9, 1.667887553E9, 1.667887601E9, 1.667887649E9, 1.667887697E9, 1.667887745E9, 1.667887793E9, 1.667887841E9, 1.667887889E9, 1.667887937E9, 1.667887985E9, 1.667888033E9, 1.667888081E9, 1.667888129E9, 1.667888177E9, 1.667888225E9, 1.667888273E9, 1.667888321E9, 1.667888369E9, 1.66788876E9, 1.667888761E9, 1.667894346E9, 1.667894394E9, 1.667894442E9, 1.66789449E9, 1.667894538E9, 1.667894586E9, 1.667894634E9, 1.667894682E9, 1.66789473E9, 1.667894778E9, 1.667894826E9, 1.667894874E9, 1.667894922E9, 1.66789497E9, 1.667895018E9, 1.667895066E9, 1.667895114E9, 1.667895162E9, 1.66789521E9, 1.667895258E9, 1.667895306E9, 1.667895354E9, 1.667895402E9, 1.66789545E9, 1.667895498E9, 1.667895546E9, 1.667895594E9, 1.667895642E9, 1.66789569E9, 1.667895738E9, 1.667895786E9, 1.667895834E9, 1.667895882E9, 1.66789593E9, 1.667895978E9, 1.667896026E9, 1.667896074E9, 1.667896122E9, 1.66789617E9, 1.667896218E9, 1.667896266E9, 1.667896314E9, 1.667896362E9, 1.66789641E9, 1.667896458E9, 1.667896506E9, 1.667896554E9, 1.667896602E9, 1.66789665E9, 1.667896698E9, 1.667896746E9, 1.667896794E9, 1.667896842E9, 1.66789689E9, 1.667896938E9, 1.667896986E9, 1.667897034E9, 1.667897082E9, 1.66789713E9, 1.667897178E9, 1.667897226E9, 1.667897274E9, 1.667897322E9, 1.66789737E9, 1.667897418E9, 1.667897466E9, 1.667897514E9, 1.667897562E9, 1.66789761E9, 1.66789794E9, 1.66789812E9, 1.667903767E9, 1.667903815E9, 1.667903863E9, 1.667903911E9, 1.667903959E9, 1.667904007E9, 1.667904055E9, 1.667904103E9, 1.667904151E9, 1.667904199E9, 1.667904247E9, 1.667904295E9, 1.667904343E9, 1.667904391E9, 1.667904439E9, 1.667904487E9, 1.667904535E9, 1.667904583E9, 1.667904631E9, 1.667904679E9, 1.667904727E9, 1.667904775E9, 1.667904823E9, 1.667904871E9, 1.667904919E9, 1.667904967E9, 1.667905015E9, 1.667905063E9, 1.667905111E9, 1.667905159E9, 1.667905207E9, 1.667905255E9, 1.667905303E9, 1.667905351E9, 1.667905399E9, 1.667905447E9, 1.667905495E9, 1.667905543E9, 1.667905591E9, 1.667905639E9, 1.667905687E9, 1.667905735E9, 1.667905783E9, 1.667905831E9, 1.667905879E9, 1.667905927E9, 1.667905975E9, 1.667906023E9, 1.667906071E9, 1.667906119E9, 1.667906167E9, 1.667906215E9, 1.667906263E9, 1.667906311E9, 1.667906359E9, 1.667906407E9, 1.667906455E9, 1.667906503E9, 1.667906551E9, 1.667906599E9, 1.667906647E9, 1.667906695E9, 1.667906743E9, 1.667906791E9, 1.667906839E9, 1.667906887E9, 1.667906935E9, 1.667906983E9, 1.667907031E9, 1.667907079E9, 1.66790736E9, 1.66790754E9, 1.667913286E9, 1.667913334E9, 1.667913382E9, 1.66791343E9, 1.667913478E9, 1.667913526E9, 1.667913574E9, 1.667913622E9, 1.66791367E9, 1.667913718E9, 1.667913766E9, 1.667913814E9, 1.667913862E9, 1.66791391E9, 1.667913958E9, 1.667914006E9, 1.667914054E9, 1.667914102E9, 1.66791415E9, 1.667914198E9, 1.667914246E9, 1.667914294E9, 1.667914342E9, 1.66791439E9, 1.667914438E9, 1.667914486E9, 1.667914534E9, 1.667914582E9, 1.66791463E9, 1.667914678E9, 1.667914726E9, 1.667914774E9, 1.667914822E9, 1.66791487E9, 1.667914918E9, 1.667914966E9, 1.667915014E9, 1.667915062E9, 1.66791511E9, 1.667915158E9, 1.667915206E9, 1.667915254E9, 1.667915302E9, 1.66791535E9, 1.667915398E9, 1.667915446E9, 1.667915494E9, 1.667915542E9, 1.66791559E9, 1.667915638E9, 1.667915686E9, 1.667915734E9, 1.667915782E9, 1.66791583E9, 1.667915878E9, 1.667915926E9, 1.667915974E9, 1.667916022E9, 1.66791607E9, 1.667916118E9, 1.667916166E9, 1.667916214E9, 1.667916262E9, 1.66791631E9, 1.667916358E9, 1.667916406E9, 1.667916454E9, 1.667916502E9, 1.66791655E9, 1.6679169E9, 1.66791714E9, 1.667923045E9, 1.667923093E9, 1.667923141E9, 1.667923189E9, 1.667923237E9, 1.667923285E9, 1.667923333E9, 1.667923381E9, 1.667923429E9, 1.667923477E9, 1.667923525E9, 1.667923573E9, 1.667923621E9, 1.667923669E9, 1.667923717E9, 1.667923765E9, 1.667923813E9, 1.667923861E9, 1.667923909E9, 1.667923957E9, 1.667924005E9, 1.667924053E9, 1.667924101E9, 1.667924149E9, 1.667924197E9, 1.667924245E9, 1.667924293E9, 1.667924341E9, 1.667924389E9, 1.667924437E9, 1.667924485E9, 1.667924533E9, 1.667924581E9, 1.667924629E9, 1.667924677E9, 1.667924725E9, 1.667924773E9, 1.667924821E9, 1.667924869E9, 1.667924917E9, 1.667924965E9, 1.667925013E9, 1.667925061E9, 1.667925109E9, 1.667925157E9, 1.667925205E9, 1.667925253E9, 1.667925301E9, 1.667925349E9, 1.667925397E9, 1.667925445E9, 1.667925493E9, 1.667925541E9, 1.667925589E9, 1.667925637E9, 1.667925685E9, 1.667925733E9, 1.667925781E9, 1.667925829E9, 1.667925877E9, 1.667925925E9, 1.667925973E9, 1.667926021E9, 1.667926069E9, 1.66792638E9, 1.66792656E9, 1.66793109E9, 1.667931138E9, 1.667931186E9, 1.667931234E9, 1.667931282E9, 1.66793133E9, 1.667931378E9, 1.667931426E9, 1.667931474E9, 1.667931522E9, 1.66793157E9, 1.667931618E9, 1.667931666E9, 1.667931714E9, 1.667931762E9, 1.66793181E9, 1.667931858E9, 1.667931906E9, 1.667931954E9, 1.667932002E9, 1.66793205E9, 1.667932098E9, 1.667932146E9, 1.667932194E9, 1.667932242E9, 1.66793229E9, 1.667932338E9, 1.667932386E9, 1.667932434E9, 1.667932482E9, 1.66793253E9, 1.667932578E9, 1.667932626E9, 1.667932674E9, 1.667932722E9, 1.66793277E9, 1.667932818E9, 1.667932866E9, 1.667932914E9, 1.667932962E9, 1.66793301E9, 1.667933058E9, 1.667933106E9, 1.667933154E9, 1.667933202E9, 1.66793325E9, 1.667933298E9, 1.667933346E9, 1.667933394E9, 1.667933442E9, 1.66793349E9, 1.66793376E9, 1.66793394E9, 1.667937572E9, 1.66793762E9, 1.667937668E9, 1.667937716E9, 1.667937764E9, 1.667937812E9, 1.66793786E9, 1.667937908E9, 1.667937956E9, 1.667938004E9, 1.667938052E9, 1.6679381E9, 1.667938148E9, 1.667938196E9, 1.667938244E9, 1.667938292E9, 1.66793834E9, 1.667938388E9, 1.667938436E9, 1.667938484E9, 1.667938532E9, 1.66793858E9, 1.667938628E9, 1.667938676E9, 1.667938724E9, 1.667938772E9, 1.66793882E9, 1.667938868E9, 1.667938916E9, 1.667938964E9, 1.667939012E9, 1.66793906E9, 1.667939108E9, 1.667939156E9, 1.667939204E9, 1.667939252E9, 1.6679393E9, 1.667939348E9, 1.667939396E9, 1.667939444E9, 1.667939492E9, 1.66793954E9, 1.66793982E9, 1.66794E9, 1.66794342E9, 1.667943468E9, 1.667943516E9, 1.667943564E9, 1.667943612E9, 1.66794366E9, 1.667943708E9, 1.667943756E9, 1.667943804E9, 1.667943852E9, 1.6679439E9, 1.667943948E9, 1.667943996E9, 1.667944044E9, 1.667944092E9, 1.66794414E9, 1.667944188E9, 1.667944236E9, 1.667944284E9, 1.667944332E9, 1.66794438E9, 1.667944428E9, 1.667944476E9, 1.667944524E9, 1.667944572E9, 1.66794462E9, 1.667944668E9, 1.667944716E9, 1.667944764E9, 1.667944812E9, 1.66794486E9, 1.667944908E9, 1.667944956E9, 1.667945004E9, 1.667945052E9, 1.6679451E9, 1.66794534E9, 1.66794546E9, 1.667948221E9, 1.667948269E9, 1.667948317E9, 1.667948365E9, 1.667948413E9, 1.667948461E9, 1.667948509E9, 1.667948557E9, 1.667948605E9, 1.667948653E9, 1.667948701E9, 1.667948749E9, 1.667948797E9, 1.667948845E9, 1.667948893E9, 1.667948941E9, 1.667948989E9, 1.667949037E9, 1.667949085E9, 1.667949133E9, 1.667949181E9, 1.667949229E9, 1.667949277E9, 1.667949325E9, 1.667949373E9, 1.667949421E9, 1.667949469E9, 1.66794972E9, 1.6679499E9, 1.667952467E9, 1.667952515E9, 1.667952563E9, 1.667952611E9, 1.667952659E9, 1.667952707E9, 1.667952755E9, 1.667952803E9, 1.667952851E9, 1.667952899E9, 1.667952947E9, 1.667952995E9, 1.667953043E9, 1.667953091E9, 1.667953139E9, 1.667953187E9, 1.667953235E9, 1.667953283E9, 1.667953331E9, 1.667953379E9, 1.667953427E9, 1.667953475E9, 1.667953523E9, 1.667953571E9, 1.667953619E9, 1.66795392E9, 1.6679541E9, 1.667956755E9, 1.667956803E9, 1.667956851E9, 1.667956899E9, 1.667956947E9, 1.667956995E9, 1.667957043E9, 1.667957091E9, 1.667957139E9, 1.667957187E9, 1.667957235E9, 1.667957283E9, 1.667957331E9, 1.667957379E9, 1.667957427E9, 1.667957475E9, 1.667957523E9, 1.667957571E9, 1.667957619E9, 1.667957667E9, 1.667957715E9, 1.667957763E9, 1.667957811E9, 1.667957859E9, 1.66795812E9, 1.6679583E9, 1.66796094E9, 1.667960988E9, 1.667961036E9, 1.667961084E9, 1.667961132E9, 1.66796118E9, 1.667961228E9, 1.667961276E9, 1.667961324E9, 1.667961372E9, 1.66796142E9, 1.667961468E9, 1.667961516E9, 1.667961564E9, 1.667961612E9, 1.66796166E9, 1.667961708E9, 1.667961756E9, 1.667961804E9, 1.667961852E9, 1.6679619E9, 1.667961948E9, 1.667961996E9, 1.667962044E9, 1.667962092E9, 1.66796214E9, 1.66796244E9, 1.66796256E9, 1.667965034E9, 1.667965082E9, 1.66796513E9, 1.667965178E9, 1.667965226E9, 1.667965274E9, 1.667965322E9, 1.66796537E9, 1.667965418E9, 1.667965466E9, 1.667965514E9, 1.667965562E9, 1.66796561E9, 1.667965658E9, 1.667965706E9, 1.667965754E9, 1.667965802E9, 1.66796585E9, 1.667965898E9, 1.667965946E9, 1.667965994E9, 1.667966042E9, 1.66796609E9, 1.66796634E9, 1.66796652E9, 1.667969196E9, 1.667969244E9, 1.667969292E9, 1.66796934E9, 1.667969388E9, 1.667969436E9, 1.667969484E9, 1.667969532E9, 1.66796958E9, 1.667969628E9, 1.667969676E9, 1.667969724E9, 1.667969772E9, 1.66796982E9, 1.667969868E9, 1.667969916E9, 1.667969964E9, 1.667970012E9, 1.66797006E9, 1.667970108E9, 1.667970156E9, 1.667970204E9, 1.667970252E9, 1.6679703E9, 1.66797054E9, 1.66797072E9, 1.667973502E9, 1.66797355E9, 1.667973598E9, 1.667973646E9, 1.667973694E9, 1.667973742E9, 1.66797379E9, 1.667973838E9, 1.667973886E9, 1.667973934E9, 1.667973982E9, 1.66797403E9, 1.667974078E9, 1.667974126E9, 1.667974174E9, 1.667974222E9, 1.66797427E9, 1.667974318E9, 1.667974366E9, 1.667974414E9, 1.667974462E9, 1.66797451E9, 1.667974558E9, 1.667974606E9, 1.667974654E9, 1.667974702E9, 1.66797475E9, 1.66797504E9, 1.66797516E9, 1.667977721E9, 1.667977769E9, 1.667977817E9, 1.667977865E9, 1.667977913E9, 1.667977961E9, 1.667978009E9, 1.667978057E9, 1.667978105E9, 1.667978153E9, 1.667978201E9, 1.667978249E9, 1.667978297E9, 1.667978345E9, 1.667978393E9, 1.667978441E9, 1.667978489E9, 1.667978537E9, 1.667978585E9, 1.667978633E9, 1.667978681E9, 1.667978729E9, 1.667978777E9, 1.667978825E9, 1.667978873E9, 1.667978921E9, 1.667978969E9, 1.66797924E9, 1.66797942E9, 1.667982191E9, 1.667982239E9, 1.667982287E9, 1.667982335E9, 1.667982383E9, 1.667982431E9, 1.667982479E9, 1.667982527E9, 1.667982575E9, 1.667982623E9, 1.667982671E9, 1.667982719E9, 1.667982767E9, 1.667982815E9, 1.667982863E9, 1.667982911E9, 1.667982959E9, 1.667983007E9, 1.667983055E9, 1.667983103E9, 1.667983151E9, 1.667983199E9, 1.66798344E9, 1.66798362E9, 1.667986021E9, 1.667986069E9, 1.667986117E9, 1.667986165E9, 1.667986213E9, 1.667986261E9, 1.667986309E9, 1.667986357E9, 1.667986405E9, 1.667986453E9, 1.667986501E9, 1.667986549E9, 1.667986597E9, 1.667986645E9, 1.667986693E9, 1.667986741E9, 1.667986789E9, 1.667986837E9, 1.667986885E9, 1.667986933E9, 1.667986981E9, 1.667987029E9, 1.667987077E9, 1.667987125E9, 1.667987173E9, 1.667987221E9, 1.667987269E9, 1.66798752E9, 1.6679877E9, 1.667990291E9, 1.667990339E9, 1.667990387E9, 1.667990435E9, 1.667990483E9, 1.667990531E9, 1.667990579E9, 1.667990627E9, 1.667990675E9, 1.667990723E9, 1.667990771E9, 1.667990819E9, 1.667990867E9, 1.667990915E9, 1.667990963E9, 1.667991011E9, 1.667991059E9, 1.667991107E9, 1.667991155E9, 1.667991203E9, 1.667991251E9, 1.667991299E9, 1.66799154E9, 1.66799166E9, 1.667994144E9, 1.667994192E9, 1.66799424E9, 1.667994288E9, 1.667994336E9, 1.667994384E9, 1.667994432E9, 1.66799448E9, 1.667994528E9, 1.667994576E9, 1.667994624E9, 1.667994672E9, 1.66799472E9, 1.667994768E9, 1.667994816E9, 1.667994864E9, 1.667994912E9, 1.66799496E9, 1.667995008E9, 1.667995056E9, 1.667995104E9, 1.667995152E9, 1.6679952E9, 1.6679955E9, 1.66799568E9, 1.667997972E9, 1.66799802E9, 1.667998068E9, 1.667998116E9, 1.667998164E9, 1.667998212E9, 1.66799826E9, 1.667998308E9, 1.667998356E9, 1.667998404E9, 1.667998452E9, 1.6679985E9, 1.667998548E9, 1.667998596E9, 1.667998644E9, 1.667998692E9, 1.66799874E9, 1.667998788E9, 1.667998836E9, 1.667998884E9, 1.667998932E9, 1.66799898E9, 1.66799922E9, 1.6679994E9, 1.668002052E9, 1.6680021E9, 1.668002148E9, 1.668002196E9, 1.668002244E9, 1.668002292E9, 1.66800234E9, 1.668002388E9, 1.668002436E9, 1.668002484E9, 1.668002532E9, 1.66800258E9, 1.668002628E9, 1.668002676E9, 1.668002724E9, 1.668002772E9, 1.66800282E9, 1.668002868E9, 1.668002916E9, 1.668002964E9, 1.668003012E9, 1.66800306E9, 1.6680033E9, 1.66800354E9, 1.668003541E9, 1.668003542E9, 1.668003543E9, 1.668003544E9, 1.668003545E9, 1.668003546E9, 1.668003547E9, 1.668003548E9, 1.668003549E9, 1.66800355E9, 1.668003551E9, 1.668003552E9, 1.668003553E9, 1.668003554E9, 1.668003555E9, 1.668003556E9, 1.668003557E9, 1.668003558E9, 1.668003559E9, 1.66800356E9, 1.668003561E9, 1.668003562E9, 1.668006855E9, 1.668006856E9, 1.66800879E9, 1.668008838E9, 1.668008886E9, 1.668008934E9, 1.668008982E9, 1.66800903E9, 1.668009078E9, 1.668009126E9, 1.668009174E9, 1.668009222E9, 1.66800927E9, 1.668009318E9, 1.668009366E9, 1.668009414E9, 1.668009462E9, 1.66800951E9, 1.668009558E9, 1.668009606E9, 1.668009654E9, 1.668009702E9, 1.66800975E9, 1.66801002E9, 1.66801026E9, 1.668010261E9, 1.668010262E9, 1.668010263E9, 1.668010264E9, 1.668010265E9, 1.668010266E9, 1.668010267E9, 1.668010268E9, 1.668010269E9, 1.66801027E9, 1.668010271E9, 1.668010272E9, 1.668010273E9, 1.668010274E9, 1.668010275E9, 1.668010276E9, 1.668010277E9, 1.668010278E9, 1.668010279E9, 1.66801028E9, 1.668010281E9, 1.668013395E9, 1.668013396E9, 1.668015218E9, 1.668015266E9, 1.668015314E9, 1.668015362E9, 1.66801541E9, 1.668015458E9, 1.668015506E9, 1.668015554E9, 1.668015602E9, 1.66801565E9, 1.668015698E9, 1.668015746E9, 1.668015794E9, 1.668015842E9, 1.66801589E9, 1.668015938E9, 1.668015986E9, 1.668016034E9, 1.668016082E9, 1.66801613E9, 1.66801638E9, 1.66801656E9, 1.668016561E9, 1.668016562E9, 1.668016563E9, 1.668016564E9, 1.668016565E9, 1.668016566E9, 1.668016567E9, 1.668016568E9, 1.668016569E9, 1.66801657E9, 1.668016571E9, 1.668016572E9, 1.668016573E9, 1.668016574E9, 1.668016575E9, 1.668016576E9, 1.668016577E9, 1.668016578E9, 1.668016579E9, 1.66801658E9, 1.668016581E9, 1.668016582E9, 1.668019671E9, 1.668019672E9, 1.668021338E9, 1.668021386E9, 1.668021434E9, 1.668021482E9, 1.66802153E9, 1.668021578E9, 1.668021626E9, 1.668021674E9, 1.668021722E9, 1.66802177E9, 1.668021818E9, 1.668021866E9, 1.668021914E9, 1.668021962E9, 1.66802201E9, 1.668022058E9, 1.668022106E9, 1.668022154E9, 1.668022202E9, 1.66802225E9, 1.6680225E9, 1.66802268E9, 1.668022681E9, 1.668022682E9, 1.668022683E9, 1.668022684E9, 1.668022685E9, 1.668022686E9, 1.668022687E9, 1.668022688E9, 1.668022689E9, 1.66802269E9, 1.668022691E9, 1.668022692E9, 1.668022693E9, 1.668022694E9, 1.668022695E9, 1.668022696E9, 1.668022697E9, 1.668022698E9, 1.668022699E9, 1.6680227E9, 1.668022701E9, 1.668025893E9, 1.668025894E9, 1.668027665E9, 1.668027713E9, 1.668027761E9, 1.668027809E9, 1.668027857E9, 1.668027905E9, 1.668027953E9, 1.668028001E9, 1.668028049E9, 1.668028097E9, 1.668028145E9, 1.668028193E9, 1.668028241E9, 1.668028289E9, 1.668028337E9, 1.668028385E9, 1.668028433E9, 1.668028481E9, 1.668028529E9, 1.6680288E9, 1.66802898E9, 1.668028981E9, 1.668028982E9, 1.668028983E9, 1.668028984E9, 1.668028985E9, 1.668028986E9, 1.668028987E9, 1.668028988E9, 1.668028989E9, 1.66802899E9, 1.668028991E9, 1.668028992E9, 1.668028993E9, 1.668028994E9, 1.668028995E9, 1.668028996E9, 1.668028997E9, 1.668028998E9, 1.668028999E9, 1.66803198E9, 1.668031981E9, 1.668033796E9, 1.668033844E9, 1.668033892E9, 1.66803394E9, 1.668033988E9, 1.668034036E9, 1.668034084E9, 1.668034132E9, 1.66803418E9, 1.668034228E9, 1.668034276E9, 1.668034324E9, 1.668034372E9, 1.66803442E9, 1.668034468E9, 1.668034516E9, 1.668034564E9, 1.668034612E9, 1.66803466E9, 1.66803498E9, 1.66803522E9, 1.668035221E9, 1.668035222E9, 1.668035223E9, 1.668035224E9, 1.668035225E9, 1.668035226E9, 1.668035227E9, 1.668035228E9, 1.668035229E9, 1.66803523E9, 1.668035231E9, 1.668035232E9, 1.668035233E9, 1.668035234E9, 1.668035235E9, 1.668035236E9, 1.668035237E9, 1.668035238E9, 1.668035239E9, 1.66803524E9, 1.668038235E9, 1.668038236E9, 1.668039996E9, 1.668040044E9, 1.668040092E9, 1.66804014E9, 1.668040188E9, 1.668040236E9, 1.668040284E9, 1.668040332E9, 1.66804038E9, 1.668040428E9, 1.668040476E9, 1.668040524E9, 1.668040572E9, 1.66804062E9, 1.668040668E9, 1.668040716E9, 1.668040764E9, 1.668040812E9, 1.66804086E9, 1.6680411E9, 1.66804128E9, 1.668041281E9, 1.668041282E9, 1.668041283E9, 1.668041284E9, 1.668041285E9, 1.668041286E9, 1.668041287E9, 1.668041288E9, 1.668041289E9, 1.66804129E9, 1.668041291E9, 1.668041292E9, 1.668041293E9, 1.668041294E9, 1.668041295E9, 1.668041296E9, 1.668041297E9, 1.668041298E9, 1.66804374E9, 1.668043741E9, 1.668043742E9, 1.668043743E9, 1.668043744E9, 1.668043745E9, 1.668043746E9, 1.668043747E9, 1.668043748E9, 1.668043749E9, 1.66804375E9, 1.668043751E9, 1.668043752E9, 1.668043753E9, 1.668043754E9, 1.668043755E9, 1.668043756E9, 1.668043757E9, 1.668043758E9, 1.668043759E9, 1.6680462E9, 1.668046201E9, 1.668047514E9, 1.668047562E9, 1.66804761E9, 1.668047658E9, 1.668047706E9, 1.668047754E9, 1.668047802E9, 1.66804785E9, 1.668047898E9, 1.668047946E9, 1.668047994E9, 1.668048042E9, 1.66804809E9, 1.668048138E9, 1.668048186E9, 1.668048234E9, 1.668048282E9, 1.66804833E9, 1.66804866E9, 1.66804884E9, 1.668048841E9, 1.668048842E9, 1.668048843E9, 1.668048844E9, 1.668048845E9, 1.668048846E9, 1.668048847E9, 1.668048848E9, 1.668048849E9, 1.66804885E9, 1.668048851E9, 1.668048852E9, 1.668048853E9, 1.668048854E9, 1.668048855E9, 1.668048856E9, 1.668048857E9, 1.668051292E9, 1.668051293E9, 1.668051294E9, 1.668051295E9, 1.668051296E9, 1.668051297E9, 1.668051298E9, 1.668051299E9, 1.6680513E9, 1.668051301E9, 1.668051302E9, 1.668051303E9, 1.668051304E9, 1.668051305E9, 1.668051306E9, 1.668051307E9, 1.668051308E9, 1.668051309E9, 1.66805131E9, 1.668051311E9, 1.668051312E9, 1.668054032E9, 1.668054033E9, 1.668055389E9, 1.668055437E9, 1.668055485E9, 1.668055533E9, 1.668055581E9, 1.668055629E9, 1.668055677E9, 1.668055725E9, 1.668055773E9, 1.668055821E9, 1.668055869E9, 1.668055917E9, 1.668055965E9, 1.668056013E9, 1.668056061E9, 1.668056109E9, 1.66805634E9, 1.66805652E9, 1.668056521E9, 1.668056522E9, 1.668056523E9, 1.668056524E9, 1.668056525E9, 1.668056526E9, 1.668056527E9, 1.668056528E9, 1.668056529E9, 1.66805653E9, 1.668056531E9, 1.668056532E9, 1.668056533E9, 1.668056534E9, 1.668056535E9, 1.668056536E9, 1.668056537E9, 1.668056538E9, 1.668056539E9, 1.66805918E9, 1.668059181E9, 1.668059182E9, 1.668059183E9, 1.668059184E9, 1.668059185E9, 1.668059186E9, 1.668059187E9, 1.668059188E9, 1.668059189E9, 1.66805919E9, 1.668059191E9, 1.668059192E9, 1.668059193E9, 1.668059194E9, 1.668059195E9, 1.668059196E9, 1.668059197E9, 1.668059198E9, 1.668059199E9, 1.6680592E9, 1.66806184E9, 1.668061841E9, 1.668063039E9, 1.668063087E9, 1.668063135E9, 1.668063183E9, 1.668063231E9, 1.668063279E9, 1.668063327E9, 1.668063375E9, 1.668063423E9, 1.668063471E9, 1.668063519E9, 1.668063567E9, 1.668063615E9, 1.668063663E9, 1.668063711E9, 1.668063759E9, 1.66806408E9, 1.66806432E9, 1.668064321E9, 1.668064322E9, 1.668064323E9, 1.668064324E9, 1.668064325E9, 1.668064326E9, 1.668064327E9, 1.668064328E9, 1.668064329E9, 1.66806433E9, 1.668064331E9, 1.668064332E9, 1.668064333E9, 1.668064334E9, 1.668064335E9, 1.668064336E9, 1.668064337E9, 1.668064338E9, 1.668064339E9, 1.668067001E9, 1.668067002E9, 1.668067003E9, 1.668067004E9, 1.668067005E9, 1.668067006E9, 1.668067007E9, 1.668067008E9, 1.668067009E9, 1.66806701E9, 1.668067011E9, 1.668067012E9, 1.668067013E9, 1.668067014E9, 1.668067015E9, 1.668067016E9, 1.668067017E9, 1.668067018E9, 1.668067019E9, 1.66806702E9, 1.668069541E9, 1.668069542E9, 1.668070892E9, 1.66807094E9, 1.668070988E9, 1.668071036E9, 1.668071084E9, 1.668071132E9, 1.66807118E9, 1.668071228E9, 1.668071276E9, 1.668071324E9, 1.668071372E9, 1.66807142E9, 1.668071468E9, 1.668071516E9, 1.668071564E9, 1.668071612E9, 1.66807166E9, 1.66807194E9, 1.66807212E9, 1.668072121E9, 1.668072122E9, 1.668072123E9, 1.668072124E9, 1.668072125E9, 1.668072126E9, 1.668072127E9, 1.668072128E9, 1.668072129E9, 1.66807213E9, 1.668072131E9, 1.668072132E9, 1.668072133E9, 1.668072134E9, 1.668072135E9, 1.668072136E9, 1.668072137E9, 1.668074588E9, 1.668074589E9, 1.66807459E9, 1.668074591E9, 1.668074592E9, 1.668074593E9, 1.668074594E9, 1.668074595E9, 1.668074596E9, 1.668074597E9, 1.668074598E9, 1.668074599E9, 1.6680746E9, 1.668074601E9, 1.668074602E9, 1.668074603E9, 1.668074604E9, 1.668074605E9, 1.668074606E9, 1.668077057E9, 1.668077058E9, 1.66807838E9, 1.668078428E9, 1.668078476E9, 1.668078524E9, 1.668078572E9, 1.66807862E9, 1.668078668E9, 1.668078716E9, 1.668078764E9, 1.668078812E9, 1.66807886E9, 1.668078908E9, 1.668078956E9, 1.668079004E9, 1.668079052E9, 1.6680791E9, 1.66807938E9, 1.66807962E9, 1.668079621E9, 1.668079622E9, 1.668079623E9, 1.668079624E9, 1.668079625E9, 1.668079626E9, 1.668079627E9, 1.668079628E9, 1.668079629E9, 1.66807963E9, 1.668079631E9, 1.668079632E9, 1.668079633E9, 1.668079634E9, 1.668079635E9, 1.668079636E9, 1.668082173E9, 1.668082174E9, 1.668082175E9, 1.668082176E9, 1.668082177E9, 1.668082178E9, 1.668082179E9, 1.66808218E9, 1.668082181E9, 1.668082182E9, 1.668082183E9, 1.668082184E9, 1.668082185E9, 1.668082186E9, 1.668082187E9, 1.668082188E9, 1.668082189E9, 1.668084566E9, 1.668084567E9, 1.668085824E9, 1.668085872E9, 1.66808592E9, 1.668085968E9, 1.668086016E9, 1.668086064E9, 1.668086112E9, 1.66808616E9, 1.668086208E9, 1.668086256E9, 1.668086304E9, 1.668086352E9, 1.6680864E9, 1.66808664E9, 1.66808682E9, 1.668086821E9, 1.668086822E9, 1.668086823E9, 1.668086824E9, 1.668086825E9, 1.668086826E9, 1.668086827E9, 1.668086828E9, 1.668086829E9, 1.66808683E9, 1.668086831E9, 1.668086832E9, 1.668086833E9, 1.668086834E9, 1.668086835E9, 1.668086836E9, 1.668086837E9, 1.6680892E9, 1.668089201E9, 1.668089202E9, 1.668089203E9, 1.668089204E9, 1.668089205E9, 1.668089206E9, 1.668089207E9, 1.668089208E9, 1.668089209E9, 1.66808921E9, 1.668089211E9, 1.668089212E9, 1.668089213E9, 1.668089214E9, 1.668089215E9, 1.668089216E9, 1.668089217E9, 1.668089218E9, 1.66809158E9, 1.668091581E9, 1.668092666E9, 1.668092714E9, 1.668092762E9, 1.66809281E9, 1.668092858E9, 1.668092906E9, 1.668092954E9, 1.668093002E9, 1.66809305E9, 1.668093098E9, 1.668093146E9, 1.668093194E9, 1.668093242E9, 1.66809329E9, 1.66809354E9, 1.66809372E9, 1.668093721E9, 1.668093722E9, 1.668093723E9, 1.668093724E9, 1.668093725E9, 1.668093726E9, 1.668093727E9, 1.668093728E9, 1.668093729E9, 1.66809373E9, 1.668093731E9, 1.668093732E9, 1.668093733E9, 1.668093734E9, 1.668093735E9, 1.66809592E9, 1.668095921E9, 1.668095922E9, 1.668095923E9, 1.668095924E9, 1.668095925E9, 1.668095926E9, 1.668095927E9, 1.668095928E9, 1.668095929E9, 1.66809593E9, 1.668095931E9, 1.668095932E9, 1.668095933E9, 1.668095934E9, 1.668095935E9, 1.668095936E9, 1.668095937E9, 1.668098267E9, 1.668098268E9, 1.668099466E9, 1.668099514E9, 1.668099562E9, 1.66809961E9, 1.668099658E9, 1.668099706E9, 1.668099754E9, 1.668099802E9, 1.66809985E9, 1.668099898E9, 1.668099946E9, 1.668099994E9, 1.668100042E9, 1.66810009E9, 1.66810032E9, 1.66810056E9, 1.668100561E9, 1.668100562E9, 1.668100563E9, 1.668100564E9, 1.668100565E9, 1.668100566E9, 1.668100567E9, 1.668100568E9, 1.668100569E9, 1.66810057E9, 1.668100571E9, 1.668100572E9, 1.668100573E9, 1.668100574E9, 1.668100575E9, 1.668100576E9, 1.668103016E9, 1.668103017E9, 1.668103018E9, 1.668103019E9, 1.66810302E9, 1.668103021E9, 1.668103022E9, 1.668103023E9, 1.668103024E9, 1.668103025E9, 1.668103026E9, 1.668103027E9, 1.668103028E9, 1.668103029E9, 1.66810303E9, 1.668103031E9, 1.668105165E9, 1.668105166E9, 1.668106333E9, 1.668106381E9, 1.668106429E9, 1.668106477E9, 1.668106525E9, 1.668106573E9, 1.668106621E9, 1.668106669E9, 1.668106717E9, 1.668106765E9, 1.668106813E9, 1.668106861E9, 1.668106909E9, 1.66810716E9, 1.66810746E9, 1.668107461E9, 1.668107462E9, 1.668107463E9, 1.668107464E9, 1.668107465E9, 1.668107466E9, 1.668107467E9, 1.668107468E9, 1.668107469E9, 1.66810747E9, 1.668107471E9, 1.668107472E9, 1.668107473E9, 1.668107474E9, 1.668107475E9, 1.668107476E9, 1.668107477E9, 1.66810984E9, 1.668109841E9, 1.668109842E9, 1.668109843E9, 1.668109844E9, 1.668109845E9, 1.668109846E9, 1.668109847E9, 1.668109848E9, 1.668109849E9, 1.66810985E9, 1.668109851E9, 1.668109852E9, 1.668109853E9, 1.668109854E9, 1.668109855E9, 1.668109856E9, 1.66811194E9, 1.668111941E9, 1.668112954E9, 1.668113002E9, 1.66811305E9, 1.668113098E9, 1.668113146E9, 1.668113194E9, 1.668113242E9, 1.66811329E9, 1.668113338E9, 1.668113386E9, 1.668113434E9, 1.668113482E9, 1.66811353E9, 1.66811376E9, 1.668114E9, 1.668114001E9, 1.668114002E9, 1.668114003E9, 1.668114004E9, 1.668114005E9, 1.668114006E9, 1.668114007E9, 1.668114008E9, 1.668114009E9, 1.66811401E9, 1.668114011E9, 1.668114012E9, 1.668114013E9, 1.668114014E9, 1.66811602E9, 1.668116021E9, 1.668116022E9, 1.668116023E9, 1.668116024E9, 1.668116025E9, 1.668116026E9, 1.668116027E9, 1.668116028E9, 1.668116029E9, 1.66811603E9, 1.668116031E9, 1.668116032E9, 1.668116033E9, 1.668116034E9, 1.668116035E9, 1.668116036E9, 1.668118184E9, 1.668118185E9, 1.668119264E9, 1.668119312E9, 1.66811936E9, 1.668119408E9, 1.668119456E9, 1.668119504E9, 1.668119552E9, 1.6681196E9, 1.668119648E9, 1.668119696E9, 1.668119744E9, 1.668119792E9, 1.66811984E9, 1.66812006E9, 1.66812042E9, 1.668120421E9, 1.668120422E9, 1.668120423E9, 1.668120424E9, 1.668120425E9, 1.668120426E9, 1.668120427E9, 1.668120428E9, 1.668120429E9, 1.66812043E9, 1.668120431E9, 1.668120432E9, 1.668120433E9, 1.66812242E9, 1.668122421E9, 1.668122422E9, 1.668122423E9, 1.668122424E9, 1.668122425E9, 1.668122426E9, 1.668122427E9, 1.668122428E9, 1.668122429E9, 1.66812243E9, 1.668122431E9, 1.668122432E9, 1.668122433E9, 1.668122434E9, 1.668122435E9, 1.668122436E9, 1.668124728E9, 1.668124729E9, 1.66812572E9, 1.668125768E9, 1.668125816E9, 1.668125864E9, 1.668125912E9, 1.66812596E9, 1.668126008E9, 1.668126056E9, 1.668126104E9, 1.668126152E9, 1.6681262E9, 1.66812642E9, 1.66812666E9, 1.668126661E9, 1.668126662E9, 1.668126663E9, 1.668126664E9, 1.668126665E9, 1.668126666E9, 1.668126667E9, 1.668126668E9, 1.668126669E9, 1.66812667E9, 1.668126671E9, 1.668126672E9, 1.668126673E9, 1.668128639E9, 1.66812864E9, 1.668128641E9, 1.668128642E9, 1.668128643E9, 1.668128644E9, 1.668128645E9, 1.668128646E9, 1.668128647E9, 1.668128648E9, 1.668128649E9, 1.66812865E9, 1.668128651E9, 1.668128652E9, 1.668128653E9, 1.668130617E9, 1.668130618E9, 1.668131958E9, 1.668132006E9, 1.668132054E9, 1.668132102E9, 1.66813215E9, 1.668132198E9, 1.668132246E9, 1.668132294E9, 1.668132342E9, 1.66813239E9, 1.668132438E9, 1.668132486E9, 1.668132534E9, 1.668132582E9, 1.66813263E9, 1.6681329E9, 1.66813308E9, 1.668133081E9, 1.668133082E9, 1.668133083E9, 1.668133084E9, 1.668133085E9, 1.668133086E9, 1.668133087E9, 1.668133088E9, 1.668133089E9, 1.66813309E9, 1.668133091E9, 1.668133092E9, 1.668133093E9, 1.668133094E9, 1.6681351E9, 1.668135101E9, 1.668135102E9, 1.668135103E9, 1.668135104E9, 1.668135105E9, 1.668135106E9, 1.668135107E9, 1.668135108E9, 1.668135109E9, 1.66813511E9, 1.668135111E9, 1.668135112E9, 1.668135113E9, 1.668135114E9, 1.668135115E9, 1.668135116E9, 1.668137264E9, 1.668137265E9, 1.668138314E9, 1.668138362E9, 1.66813841E9, 1.668138458E9, 1.668138506E9, 1.668138554E9, 1.668138602E9, 1.66813865E9, 1.668138698E9, 1.668138746E9, 1.668138794E9, 1.668138842E9, 1.66813889E9, 1.66813914E9, 1.66813938E9, 1.668139381E9, 1.668139382E9, 1.668139383E9, 1.668139384E9, 1.668139385E9, 1.668139386E9, 1.668139387E9, 1.668139388E9, 1.668139389E9, 1.66813939E9, 1.668139391E9, 1.668139392E9, 1.668139393E9, 1.668139394E9, 1.66814148E9, 1.668141481E9, 1.668141482E9, 1.668141483E9, 1.668141484E9, 1.668141485E9, 1.668141486E9, 1.668141487E9, 1.668141488E9, 1.668141489E9, 1.66814149E9, 1.668141491E9, 1.668141492E9, 1.668141493E9, 1.668141494E9, 1.668141495E9, 1.66814358E9, 1.668143581E9, 1.668144806E9, 1.668144854E9, 1.668144902E9, 1.66814495E9, 1.668144998E9, 1.668145046E9, 1.668145094E9, 1.668145142E9, 1.66814519E9, 1.668145238E9, 1.668145286E9, 1.668145334E9, 1.668145382E9, 1.66814543E9, 1.66814568E9, 1.66814604E9, 1.668146041E9, 1.668146042E9, 1.668146043E9, 1.668146044E9, 1.668146045E9, 1.668146046E9, 1.668146047E9, 1.668146048E9, 1.668146049E9, 1.66814605E9, 1.668146051E9, 1.668146052E9, 1.668146053E9, 1.668146054E9, 1.668146055E9, 1.668146056E9, 1.66814838E9, 1.668148381E9, 1.668148382E9, 1.668148383E9, 1.668148384E9, 1.668148385E9, 1.668148386E9, 1.668148387E9, 1.668148388E9, 1.668148389E9, 1.66814839E9, 1.668148391E9, 1.668148392E9, 1.668148393E9, 1.668148394E9, 1.668148395E9, 1.668148396E9, 1.668148397E9, 1.66815072E9, 1.668150721E9, 1.668152059E9, 1.668152107E9, 1.668152155E9, 1.668152203E9, 1.668152251E9, 1.668152299E9, 1.668152347E9, 1.668152395E9, 1.668152443E9, 1.668152491E9, 1.668152539E9, 1.668152587E9, 1.668152635E9, 1.668152683E9, 1.668152731E9, 1.668152779E9, 1.66815306E9, 1.6681533E9, 1.668153301E9, 1.668153302E9, 1.668153303E9, 1.668153304E9, 1.668153305E9, 1.668153306E9, 1.668153307E9, 1.668153308E9, 1.668153309E9, 1.66815331E9, 1.668153311E9, 1.668153312E9, 1.668153313E9, 1.668153314E9, 1.668153315E9, 1.668153316E9, 1.668153317E9, 1.66815583E9, 1.668155831E9, 1.668155832E9, 1.668155833E9, 1.668155834E9, 1.668155835E9, 1.668155836E9, 1.668155837E9, 1.668155838E9, 1.668155839E9, 1.66815584E9, 1.668155841E9, 1.668155842E9, 1.668155843E9, 1.668155844E9, 1.668155845E9, 1.668155846E9, 1.668155847E9, 1.668155848E9, 1.668158359E9, 1.66815836E9, 1.66815973E9, 1.668159778E9, 1.668159826E9, 1.668159874E9, 1.668159922E9, 1.66815997E9, 1.668160018E9, 1.668160066E9, 1.668160114E9, 1.668160162E9, 1.66816021E9, 1.668160258E9, 1.668160306E9, 1.668160354E9, 1.668160402E9, 1.66816045E9, 1.66816074E9, 1.66816092E9, 1.668160921E9, 1.668160922E9, 1.668160923E9, 1.668160924E9, 1.668160925E9, 1.668160926E9, 1.668160927E9, 1.668160928E9, 1.668160929E9, 1.66816093E9, 1.668160931E9, 1.668160932E9, 1.668160933E9, 1.668160934E9, 1.668160935E9, 1.668160936E9, 1.668160937E9, 1.668160938E9, 1.668163599E9, 1.6681636E9, 1.668163601E9, 1.668163602E9, 1.668163603E9, 1.668163604E9, 1.668163605E9, 1.668163606E9, 1.668163607E9, 1.668163608E9, 1.668163609E9, 1.66816361E9, 1.668163611E9, 1.668163612E9, 1.668163613E9, 1.668163614E9, 1.668163615E9, 1.668163616E9, 1.668163617E9, 1.668163618E9, 1.668166278E9, 1.668166279E9, 1.6681676E9, 1.668167648E9, 1.668167696E9, 1.668167744E9, 1.668167792E9, 1.66816784E9, 1.668167888E9, 1.668167936E9, 1.668167984E9, 1.668168032E9, 1.66816808E9, 1.668168128E9, 1.668168176E9, 1.668168224E9, 1.668168272E9, 1.66816832E9, 1.66816866E9, 1.6681689E9, 1.668168901E9, 1.668168902E9, 1.668168903E9, 1.668168904E9, 1.668168905E9, 1.668168906E9, 1.668168907E9, 1.668168908E9, 1.668168909E9, 1.66816891E9, 1.668168911E9, 1.668168912E9, 1.668168913E9, 1.668168914E9, 1.668168915E9, 1.668168916E9, 1.668168917E9, 1.668168918E9, 1.668168919E9, 1.668171534E9, 1.668171535E9, 1.668171536E9, 1.668171537E9, 1.668171538E9, 1.668171539E9, 1.66817154E9, 1.668171541E9, 1.668171542E9, 1.668171543E9, 1.668171544E9, 1.668171545E9, 1.668171546E9, 1.668171547E9, 1.668171548E9, 1.668171549E9, 1.66817155E9, 1.668171551E9, 1.668171552E9, 1.668171553E9, 1.668171554E9, 1.668174168E9, 1.668174169E9, 1.668175758E9, 1.668175806E9, 1.668175854E9, 1.668175902E9, 1.66817595E9, 1.668175998E9, 1.668176046E9, 1.668176094E9, 1.668176142E9, 1.66817619E9, 1.668176238E9, 1.668176286E9, 1.668176334E9, 1.668176382E9, 1.66817643E9, 1.668176478E9, 1.668176526E9, 1.668176574E9, 1.668176622E9, 1.66817667E9, 1.66817694E9, 1.66817724E9, 1.668177241E9, 1.668177242E9, 1.668177243E9, 1.668177244E9, 1.668177245E9, 1.668177246E9, 1.668177247E9, 1.668177248E9, 1.668177249E9, 1.66817725E9, 1.668177251E9, 1.668177252E9, 1.668177253E9, 1.668177254E9, 1.668177255E9, 1.668177256E9, 1.668177257E9, 1.668177258E9, 1.668177259E9, 1.66817726E9, 1.668177261E9, 1.668180296E9, 1.668180297E9, 1.668181945E9, 1.668181993E9, 1.668182041E9, 1.668182089E9, 1.668182137E9, 1.668182185E9, 1.668182233E9, 1.668182281E9, 1.668182329E9, 1.668182377E9, 1.668182425E9, 1.668182473E9, 1.668182521E9, 1.668182569E9, 1.668182617E9, 1.668182665E9, 1.668182713E9, 1.668182761E9, 1.668182809E9, 1.66818306E9, 1.6681833E9, 1.668183301E9, 1.668183302E9, 1.668183303E9, 1.668183304E9, 1.668183305E9, 1.668183306E9, 1.668183307E9, 1.668183308E9, 1.668183309E9, 1.66818331E9, 1.668183311E9, 1.668183312E9, 1.668183313E9, 1.668183314E9, 1.668183315E9, 1.668183316E9, 1.668183317E9, 1.668183318E9, 1.668183319E9, 1.66818332E9, 1.668183321E9, 1.668183322E9, 1.668183323E9, 1.668183324E9, 1.668186548E9, 1.668186549E9, 1.668188323E9, 1.668188371E9, 1.668188419E9, 1.668188467E9, 1.668188515E9, 1.668188563E9, 1.668188611E9, 1.668188659E9, 1.668188707E9, 1.668188755E9, 1.668188803E9, 1.668188851E9, 1.668188899E9, 1.668188947E9, 1.668188995E9, 1.668189043E9, 1.668189091E9, 1.668189139E9, 1.668189187E9, 1.668189235E9, 1.668189283E9, 1.668189331E9, 1.668189379E9, 1.66818966E9, 1.66818984E9, 1.668189841E9, 1.668189842E9, 1.668189843E9, 1.668189844E9, 1.668189845E9, 1.668189846E9, 1.668189847E9, 1.668189848E9, 1.668189849E9, 1.66818985E9, 1.668189851E9, 1.668189852E9, 1.668189853E9, 1.668189854E9, 1.668189855E9, 1.668189856E9, 1.668189857E9, 1.668189858E9, 1.668189859E9, 1.66818986E9, 1.668189861E9, 1.668189862E9, 1.668189863E9, 1.668189864E9, 1.66819326E9, 1.668193261E9, 1.668195336E9, 1.668195384E9, 1.668195432E9, 1.66819548E9, 1.668195528E9, 1.668195576E9, 1.668195624E9, 1.668195672E9, 1.66819572E9, 1.668195768E9, 1.668195816E9, 1.668195864E9, 1.668195912E9, 1.66819596E9, 1.668196008E9, 1.668196056E9, 1.668196104E9, 1.668196152E9, 1.6681962E9, 1.668196248E9, 1.668196296E9, 1.668196344E9, 1.668196392E9, 1.66819644E9, 1.66819668E9, 1.66819686E9, 1.668196861E9, 1.668196862E9, 1.668196863E9, 1.668196864E9, 1.668196865E9, 1.668196866E9, 1.668196867E9, 1.668196868E9, 1.668196869E9, 1.66819687E9, 1.668196871E9, 1.668196872E9, 1.668196873E9, 1.668196874E9, 1.668196875E9, 1.668196876E9, 1.668196877E9, 1.668196878E9, 1.668196879E9, 1.66819688E9, 1.668196881E9, 1.668196882E9, 1.668196883E9, 1.668196884E9, 1.668196885E9, 1.668196886E9, 1.66820043E9, 1.668200431E9, 1.668202549E9, 1.668202597E9, 1.668202645E9, 1.668202693E9, 1.668202741E9, 1.668202789E9, 1.668202837E9, 1.668202885E9, 1.668202933E9, 1.668202981E9, 1.668203029E9, 1.668203077E9, 1.668203125E9, 1.668203173E9, 1.668203221E9, 1.668203269E9, 1.668203317E9, 1.668203365E9, 1.668203413E9, 1.668203461E9, 1.668203509E9, 1.668203557E9, 1.668203605E9, 1.668203653E9, 1.668203701E9, 1.668203749E9, 1.668204E9, 1.668207941E9, 1.668210108E9, 1.668210156E9, 1.668210204E9, 1.668210252E9, 1.6682103E9, 1.668210348E9, 1.668210396E9, 1.668210444E9, 1.668210492E9, 1.66821054E9, 1.668210588E9, 1.668210636E9, 1.668210684E9, 1.668210732E9, 1.66821078E9, 1.668210828E9, 1.668210876E9, 1.668210924E9, 1.668210972E9, 1.66821102E9, 1.668211068E9, 1.668211116E9, 1.668211164E9, 1.668211212E9, 1.66821126E9, 1.6682115E9, 1.66821174E9, 1.668211741E9, 1.668211742E9, 1.668211743E9, 1.668211744E9, 1.668211745E9, 1.668211746E9, 1.668211747E9, 1.668211748E9, 1.668211749E9, 1.66821175E9, 1.668211751E9, 1.668211752E9, 1.668211753E9, 1.668211754E9, 1.668211755E9, 1.668211756E9, 1.668211757E9, 1.668211758E9, 1.668211759E9, 1.66821176E9, 1.668211761E9, 1.668211762E9, 1.668211763E9, 1.668211764E9, 1.668211765E9, 1.668211766E9, 1.668211767E9, 1.668215472E9, 1.668215473E9, 1.668217855E9, 1.668217903E9, 1.668217951E9, 1.668217999E9, 1.668218047E9, 1.668218095E9, 1.668218143E9, 1.668218191E9, 1.668218239E9, 1.668218287E9, 1.668218335E9, 1.668218383E9, 1.668218431E9, 1.668218479E9, 1.668218527E9, 1.668218575E9, 1.668218623E9, 1.668218671E9, 1.668218719E9, 1.668218767E9, 1.668218815E9, 1.668218863E9, 1.668218911E9, 1.668218959E9, 1.668219007E9, 1.668219055E9, 1.668219103E9, 1.668219151E9, 1.668219199E9, 1.66821948E9, 1.66821972E9, 1.668219721E9, 1.668219722E9, 1.668219723E9, 1.668219724E9, 1.668219725E9, 1.668219726E9, 1.668219727E9, 1.668219728E9, 1.668219729E9, 1.66821973E9, 1.668219731E9, 1.668219732E9, 1.668219733E9, 1.668219734E9, 1.668219735E9, 1.668219736E9, 1.668219737E9, 1.668219738E9, 1.668219739E9, 1.66821974E9, 1.668219741E9, 1.668219742E9, 1.668219743E9, 1.668219744E9, 1.668219745E9, 1.668219746E9, 1.668219747E9, 1.668219748E9, 1.668219749E9, 1.66821975E9, 1.668219751E9, 1.668219752E9, 1.668219753E9, 1.668219754E9, 1.668224297E9, 1.668224298E9, 1.668227916E9, 1.668227964E9, 1.668228012E9, 1.66822806E9, 1.668228108E9, 1.668228156E9, 1.668228204E9, 1.668228252E9, 1.6682283E9, 1.668228348E9, 1.668228396E9, 1.668228444E9, 1.668228492E9, 1.66822854E9, 1.668228588E9, 1.668228636E9, 1.668228684E9, 1.668228732E9, 1.66822878E9, 1.668228828E9, 1.668228876E9, 1.668228924E9, 1.668228972E9, 1.66822902E9, 1.668229068E9, 1.668229116E9, 1.668229164E9, 1.668229212E9, 1.66822926E9, 1.668229308E9, 1.668229356E9, 1.668229404E9, 1.668229452E9, 1.6682295E9, 1.668229548E9, 1.668229596E9, 1.668229644E9, 1.668229692E9, 1.66822974E9, 1.668229788E9, 1.668229836E9, 1.668229884E9, 1.668229932E9, 1.66822998E9, 1.66823022E9, 1.6682304E9, 1.668235263E9, 1.668235311E9, 1.668235359E9, 1.668235407E9, 1.668235455E9, 1.668235503E9, 1.668235551E9, 1.668235599E9, 1.668235647E9, 1.668235695E9, 1.668235743E9, 1.668235791E9, 1.668235839E9, 1.668235887E9, 1.668235935E9, 1.668235983E9, 1.668236031E9, 1.668236079E9, 1.668236127E9, 1.668236175E9, 1.668236223E9, 1.668236271E9, 1.668236319E9, 1.668236367E9, 1.668236415E9, 1.668236463E9, 1.668236511E9, 1.668236559E9, 1.668236607E9, 1.668236655E9, 1.668236703E9, 1.668236751E9, 1.668236799E9, 1.668236847E9, 1.668236895E9, 1.668236943E9, 1.668236991E9, 1.668237039E9, 1.668237087E9, 1.668237135E9, 1.668237183E9, 1.668237231E9, 1.668237279E9, 1.668237327E9, 1.668237375E9, 1.668237423E9, 1.668237471E9, 1.668237519E9, 1.668237567E9, 1.668237615E9, 1.668237663E9, 1.668237711E9, 1.668237759E9, 1.66823808E9, 1.66823826E9, 1.668243683E9, 1.668243731E9, 1.668243779E9, 1.668243827E9, 1.668243875E9, 1.668243923E9, 1.668243971E9, 1.668244019E9, 1.668244067E9, 1.668244115E9, 1.668244163E9, 1.668244211E9, 1.668244259E9, 1.668244307E9, 1.668244355E9, 1.668244403E9, 1.668244451E9, 1.668244499E9, 1.668244547E9, 1.668244595E9, 1.668244643E9, 1.668244691E9, 1.668244739E9, 1.668244787E9, 1.668244835E9, 1.668244883E9, 1.668244931E9, 1.668244979E9, 1.668245027E9, 1.668245075E9, 1.668245123E9, 1.668245171E9, 1.668245219E9, 1.668245267E9, 1.668245315E9, 1.668245363E9, 1.668245411E9, 1.668245459E9, 1.668245507E9, 1.668245555E9, 1.668245603E9, 1.668245651E9, 1.668245699E9, 1.668245747E9, 1.668245795E9, 1.668245843E9, 1.668245891E9, 1.668245939E9, 1.668245987E9, 1.668246035E9, 1.668246083E9, 1.668246131E9, 1.668246179E9, 1.668246227E9, 1.668246275E9, 1.668246323E9, 1.668246371E9, 1.668246419E9, 1.668246467E9, 1.668246515E9, 1.668246563E9, 1.668246611E9, 1.668246659E9, 1.668246707E9, 1.668246755E9, 1.668246803E9, 1.668246851E9, 1.668246899E9, 1.66824732E9, 1.6682475E9, 1.668253324E9, 1.668253372E9, 1.66825342E9, 1.668253468E9, 1.668253516E9, 1.668253564E9, 1.668253612E9, 1.66825366E9, 1.668253708E9, 1.668253756E9, 1.668253804E9, 1.668253852E9, 1.6682539E9, 1.668253948E9, 1.668253996E9, 1.668254044E9, 1.668254092E9, 1.66825414E9, 1.668254188E9, 1.668254236E9, 1.668254284E9, 1.668254332E9, 1.66825438E9, 1.668254428E9, 1.668254476E9, 1.668254524E9, 1.668254572E9, 1.66825462E9, 1.668254668E9, 1.668254716E9, 1.668254764E9, 1.668254812E9, 1.66825486E9, 1.668254908E9, 1.668254956E9, 1.668255004E9, 1.668255052E9, 1.6682551E9, 1.668255148E9, 1.668255196E9, 1.668255244E9, 1.668255292E9, 1.66825534E9, 1.668255388E9, 1.668255436E9, 1.668255484E9, 1.668255532E9, 1.66825558E9, 1.668255628E9, 1.668255676E9, 1.668255724E9, 1.668255772E9, 1.66825582E9, 1.668255868E9, 1.668255916E9, 1.668255964E9, 1.668256012E9, 1.66825606E9, 1.668256108E9, 1.668256156E9, 1.668256204E9, 1.668256252E9, 1.6682563E9, 1.668256348E9, 1.668256396E9, 1.668256444E9, 1.668256492E9, 1.66825654E9, 1.66825686E9, 1.6682571E9, 1.668262632E9, 1.66826268E9, 1.668262728E9, 1.668262776E9, 1.668262824E9, 1.668262872E9, 1.66826292E9, 1.668262968E9, 1.668263016E9, 1.668263064E9, 1.668263112E9, 1.66826316E9, 1.668263208E9, 1.668263256E9, 1.668263304E9, 1.668263352E9, 1.6682634E9, 1.668263448E9, 1.668263496E9, 1.668263544E9, 1.668263592E9, 1.66826364E9, 1.668263688E9, 1.668263736E9, 1.668263784E9, 1.668263832E9, 1.66826388E9, 1.668263928E9, 1.668263976E9, 1.668264024E9, 1.668264072E9, 1.66826412E9, 1.668264168E9, 1.668264216E9, 1.668264264E9, 1.668264312E9, 1.66826436E9, 1.668264408E9, 1.668264456E9, 1.668264504E9, 1.668264552E9, 1.6682646E9, 1.668264648E9, 1.668264696E9, 1.668264744E9, 1.668264792E9, 1.66826484E9, 1.668264888E9, 1.668264936E9, 1.668264984E9, 1.668265032E9, 1.66826508E9, 1.668265128E9, 1.668265176E9, 1.668265224E9, 1.668265272E9, 1.66826532E9, 1.668265368E9, 1.668265416E9, 1.668265464E9, 1.668265512E9, 1.66826556E9, 1.668265608E9, 1.668265656E9, 1.668265704E9, 1.668265752E9, 1.6682658E9, 1.66826616E9, 1.66826646E9, 1.668272312E9, 1.66827236E9, 1.668272408E9, 1.668272456E9, 1.668272504E9, 1.668272552E9, 1.6682726E9, 1.668272648E9, 1.668272696E9, 1.668272744E9, 1.668272792E9, 1.66827284E9, 1.668272888E9, 1.668272936E9, 1.668272984E9, 1.668273032E9, 1.66827308E9, 1.668273128E9, 1.668273176E9, 1.668273224E9, 1.668273272E9, 1.66827332E9, 1.668273368E9, 1.668273416E9, 1.668273464E9, 1.668273512E9, 1.66827356E9, 1.668273608E9, 1.668273656E9, 1.668273704E9, 1.668273752E9, 1.6682738E9, 1.668273848E9, 1.668273896E9, 1.668273944E9, 1.668273992E9, 1.66827404E9, 1.668274088E9, 1.668274136E9, 1.668274184E9, 1.668274232E9, 1.66827428E9, 1.668274328E9, 1.668274376E9, 1.668274424E9, 1.668274472E9, 1.66827452E9, 1.668274568E9, 1.668274616E9, 1.668274664E9, 1.668274712E9, 1.66827476E9, 1.668274808E9, 1.668274856E9, 1.668274904E9, 1.668274952E9, 1.668275E9, 1.668275048E9, 1.668275096E9, 1.668275144E9, 1.668275192E9, 1.66827524E9, 1.668275288E9, 1.668275336E9, 1.668275384E9, 1.668275432E9, 1.66827548E9, 1.66827582E9, 1.66827606E9, 1.668281665E9, 1.668281713E9, 1.668281761E9, 1.668281809E9, 1.668281857E9, 1.668281905E9, 1.668281953E9, 1.668282001E9, 1.668282049E9, 1.668282097E9, 1.668282145E9, 1.668282193E9, 1.668282241E9, 1.668282289E9, 1.668282337E9, 1.668282385E9, 1.668282433E9, 1.668282481E9, 1.668282529E9, 1.668282577E9, 1.668282625E9, 1.668282673E9, 1.668282721E9, 1.668282769E9, 1.668282817E9, 1.668282865E9, 1.668282913E9, 1.668282961E9, 1.668283009E9, 1.668283057E9, 1.668283105E9, 1.668283153E9, 1.668283201E9, 1.668283249E9, 1.668283297E9, 1.668283345E9, 1.668283393E9, 1.668283441E9, 1.668283489E9, 1.668283537E9, 1.668283585E9, 1.668283633E9, 1.668283681E9, 1.668283729E9, 1.668283777E9, 1.668283825E9, 1.668283873E9, 1.668283921E9, 1.668283969E9, 1.668284017E9, 1.668284065E9, 1.668284113E9, 1.668284161E9, 1.668284209E9, 1.668284257E9, 1.668284305E9, 1.668284353E9, 1.668284401E9, 1.668284449E9, 1.668284497E9, 1.668284545E9, 1.668284593E9, 1.668284641E9, 1.668284689E9, 1.668284737E9, 1.668284785E9, 1.668284833E9, 1.668284881E9, 1.668284929E9, 1.6682853E9, 1.66828548E9, 1.668291271E9, 1.668291319E9, 1.668291367E9, 1.668291415E9, 1.668291463E9, 1.668291511E9, 1.668291559E9, 1.668291607E9, 1.668291655E9, 1.668291703E9, 1.668291751E9, 1.668291799E9, 1.668291847E9, 1.668291895E9, 1.668291943E9, 1.668291991E9, 1.668292039E9, 1.668292087E9, 1.668292135E9, 1.668292183E9, 1.668292231E9, 1.668292279E9, 1.668292327E9, 1.668292375E9, 1.668292423E9, 1.668292471E9, 1.668292519E9, 1.668292567E9, 1.668292615E9, 1.668292663E9, 1.668292711E9, 1.668292759E9, 1.668292807E9, 1.668292855E9, 1.668292903E9, 1.668292951E9, 1.668292999E9, 1.668293047E9, 1.668293095E9, 1.668293143E9, 1.668293191E9, 1.668293239E9, 1.668293287E9, 1.668293335E9, 1.668293383E9, 1.668293431E9, 1.668293479E9, 1.668293527E9, 1.668293575E9, 1.668293623E9, 1.668293671E9, 1.668293719E9, 1.668293767E9, 1.668293815E9, 1.668293863E9, 1.668293911E9, 1.668293959E9, 1.668294007E9, 1.668294055E9, 1.668294103E9, 1.668294151E9, 1.668294199E9, 1.668294247E9, 1.668294295E9, 1.668294343E9, 1.668294391E9, 1.668294439E9, 1.66829478E9, 1.66829496E9, 1.668300898E9, 1.668300946E9, 1.668300994E9, 1.668301042E9, 1.66830109E9, 1.668301138E9, 1.668301186E9, 1.668301234E9, 1.668301282E9, 1.66830133E9, 1.668301378E9, 1.668301426E9, 1.668301474E9, 1.668301522E9, 1.66830157E9, 1.668301618E9, 1.668301666E9, 1.668301714E9, 1.668301762E9, 1.66830181E9, 1.668301858E9, 1.668301906E9, 1.668301954E9, 1.668302002E9, 1.66830205E9, 1.668302098E9, 1.668302146E9, 1.668302194E9, 1.668302242E9, 1.66830229E9, 1.668302338E9, 1.668302386E9, 1.668302434E9, 1.668302482E9, 1.66830253E9, 1.668302578E9, 1.668302626E9, 1.668302674E9, 1.668302722E9, 1.66830277E9, 1.668302818E9, 1.668302866E9, 1.668302914E9, 1.668302962E9, 1.66830301E9, 1.668303058E9, 1.668303106E9, 1.668303154E9, 1.668303202E9, 1.66830325E9, 1.668303298E9, 1.668303346E9, 1.668303394E9, 1.668303442E9, 1.66830349E9, 1.668303538E9, 1.668303586E9, 1.668303634E9, 1.668303682E9, 1.66830373E9, 1.668303778E9, 1.668303826E9, 1.668303874E9, 1.668303922E9, 1.66830397E9, 1.668304018E9, 1.668304066E9, 1.668304114E9, 1.668304162E9, 1.66830421E9, 1.6683045E9, 1.66830468E9, 1.668310557E9, 1.668310605E9, 1.668310653E9, 1.668310701E9, 1.668310749E9, 1.668310797E9, 1.668310845E9, 1.668310893E9, 1.668310941E9, 1.668310989E9, 1.668311037E9, 1.668311085E9, 1.668311133E9, 1.668311181E9, 1.668311229E9, 1.668311277E9, 1.668311325E9, 1.668311373E9, 1.668311421E9, 1.668311469E9, 1.668311517E9, 1.668311565E9, 1.668311613E9, 1.668311661E9, 1.668311709E9, 1.668311757E9, 1.668311805E9, 1.668311853E9, 1.668311901E9, 1.668311949E9, 1.668311997E9, 1.668312045E9, 1.668312093E9, 1.668312141E9, 1.668312189E9, 1.668312237E9, 1.668312285E9, 1.668312333E9, 1.668312381E9, 1.668312429E9, 1.668312477E9, 1.668312525E9, 1.668312573E9, 1.668312621E9, 1.668312669E9, 1.668312717E9, 1.668312765E9, 1.668312813E9, 1.668312861E9, 1.668312909E9, 1.668312957E9, 1.668313005E9, 1.668313053E9, 1.668313101E9, 1.668313149E9, 1.668313197E9, 1.668313245E9, 1.668313293E9, 1.668313341E9, 1.668313389E9, 1.668313437E9, 1.668313485E9, 1.668313533E9, 1.668313581E9, 1.668313629E9, 1.66831398E9, 1.66831416E9, 1.668319951E9, 1.668319999E9, 1.668320047E9, 1.668320095E9, 1.668320143E9, 1.668320191E9, 1.668320239E9, 1.668320287E9, 1.668320335E9, 1.668320383E9, 1.668320431E9, 1.668320479E9, 1.668320527E9, 1.668320575E9, 1.668320623E9, 1.668320671E9, 1.668320719E9, 1.668320767E9, 1.668320815E9, 1.668320863E9, 1.668320911E9, 1.668320959E9, 1.668321007E9, 1.668321055E9, 1.668321103E9, 1.668321151E9, 1.668321199E9, 1.668321247E9, 1.668321295E9, 1.668321343E9, 1.668321391E9, 1.668321439E9, 1.668321487E9, 1.668321535E9, 1.668321583E9, 1.668321631E9, 1.668321679E9, 1.668321727E9, 1.668321775E9, 1.668321823E9, 1.668321871E9, 1.668321919E9, 1.668321967E9, 1.668322015E9, 1.668322063E9, 1.668322111E9, 1.668322159E9, 1.668322207E9, 1.668322255E9, 1.668322303E9, 1.668322351E9, 1.668322399E9, 1.668322447E9, 1.668322495E9, 1.668322543E9, 1.668322591E9, 1.668322639E9, 1.668322687E9, 1.668322735E9, 1.668322783E9, 1.668322831E9, 1.668322879E9, 1.668322927E9, 1.668322975E9, 1.668323023E9, 1.668323071E9, 1.668323119E9, 1.66832346E9, 1.66832364E9, 1.668329317E9, 1.668329365E9, 1.668329413E9, 1.668329461E9, 1.668329509E9, 1.668329557E9, 1.668329605E9, 1.668329653E9, 1.668329701E9, 1.668329749E9, 1.668329797E9, 1.668329845E9, 1.668329893E9, 1.668329941E9, 1.668329989E9, 1.668330037E9, 1.668330085E9, 1.668330133E9, 1.668330181E9, 1.668330229E9, 1.668330277E9, 1.668330325E9, 1.668330373E9, 1.668330421E9, 1.668330469E9, 1.668330517E9, 1.668330565E9, 1.668330613E9, 1.668330661E9, 1.668330709E9, 1.668330757E9, 1.668330805E9, 1.668330853E9, 1.668330901E9, 1.668330949E9, 1.668330997E9, 1.668331045E9, 1.668331093E9, 1.668331141E9, 1.668331189E9, 1.668331237E9, 1.668331285E9, 1.668331333E9, 1.668331381E9, 1.668331429E9, 1.668331477E9, 1.668331525E9, 1.668331573E9, 1.668331621E9, 1.668331669E9, 1.668331717E9, 1.668331765E9, 1.668331813E9, 1.668331861E9, 1.668331909E9, 1.668331957E9, 1.668332005E9, 1.668332053E9, 1.668332101E9, 1.668332149E9, 1.668332197E9, 1.668332245E9, 1.668332293E9, 1.668332341E9, 1.668332389E9, 1.668332437E9, 1.668332485E9, 1.668332533E9, 1.668332581E9, 1.668332629E9, 1.66833294E9, 1.66833312E9, 1.6683386E9, 1.668338648E9, 1.668338696E9, 1.668338744E9, 1.668338792E9, 1.66833884E9, 1.668338888E9, 1.668338936E9, 1.668338984E9, 1.668339032E9, 1.66833908E9, 1.668339128E9, 1.668339176E9, 1.668339224E9, 1.668339272E9, 1.66833932E9, 1.668339368E9, 1.668339416E9, 1.668339464E9, 1.668339512E9, 1.66833956E9, 1.668339608E9, 1.668339656E9, 1.668339704E9, 1.668339752E9, 1.6683398E9, 1.668339848E9, 1.668339896E9, 1.668339944E9, 1.668339992E9, 1.66834004E9, 1.668340088E9, 1.668340136E9, 1.668340184E9, 1.668340232E9, 1.66834028E9, 1.668340328E9, 1.668340376E9, 1.668340424E9, 1.668340472E9, 1.66834052E9, 1.668340568E9, 1.668340616E9, 1.668340664E9, 1.668340712E9, 1.66834076E9, 1.668340808E9, 1.668340856E9, 1.668340904E9, 1.668340952E9, 1.668341E9, 1.668341048E9, 1.668341096E9, 1.668341144E9, 1.668341192E9, 1.66834124E9, 1.668341288E9, 1.668341336E9, 1.668341384E9, 1.668341432E9, 1.66834148E9, 1.668341528E9, 1.668341576E9, 1.668341624E9, 1.668341672E9, 1.66834172E9, 1.668341768E9, 1.668341816E9, 1.668341864E9, 1.668341912E9, 1.66834196E9, 1.6683423E9, 1.66834248E9, 1.668348054E9, 1.668348102E9, 1.66834815E9, 1.668348198E9, 1.668348246E9, 1.668348294E9, 1.668348342E9, 1.66834839E9, 1.668348438E9, 1.668348486E9, 1.668348534E9, 1.668348582E9, 1.66834863E9, 1.668348678E9, 1.668348726E9, 1.668348774E9, 1.668348822E9, 1.66834887E9, 1.668348918E9, 1.668348966E9, 1.668349014E9, 1.668349062E9, 1.66834911E9, 1.668349158E9, 1.668349206E9, 1.668349254E9, 1.668349302E9, 1.66834935E9, 1.668349398E9, 1.668349446E9, 1.668349494E9, 1.668349542E9, 1.66834959E9, 1.668349638E9, 1.668349686E9, 1.668349734E9, 1.668349782E9, 1.66834983E9, 1.668349878E9, 1.668349926E9, 1.668349974E9, 1.668350022E9, 1.66835007E9, 1.668350118E9, 1.668350166E9, 1.668350214E9, 1.668350262E9, 1.66835031E9, 1.668350358E9, 1.668350406E9, 1.668350454E9, 1.668350502E9, 1.66835055E9, 1.668350598E9, 1.668350646E9, 1.668350694E9, 1.668350742E9, 1.66835079E9, 1.668350838E9, 1.668350886E9, 1.668350934E9, 1.668350982E9, 1.66835103E9, 1.668351078E9, 1.668351126E9, 1.668351174E9, 1.668351222E9, 1.66835127E9, 1.6683516E9, 1.66835172E9, 1.668357553E9, 1.668357601E9, 1.668357649E9, 1.668357697E9, 1.668357745E9, 1.668357793E9, 1.668357841E9, 1.668357889E9, 1.668357937E9, 1.668357985E9, 1.668358033E9, 1.668358081E9, 1.668358129E9, 1.668358177E9, 1.668358225E9, 1.668358273E9, 1.668358321E9, 1.668358369E9, 1.668358417E9, 1.668358465E9, 1.668358513E9, 1.668358561E9, 1.668358609E9, 1.668358657E9, 1.668358705E9, 1.668358753E9, 1.668358801E9, 1.668358849E9, 1.668358897E9, 1.668358945E9, 1.668358993E9, 1.668359041E9, 1.668359089E9, 1.668359137E9, 1.668359185E9, 1.668359233E9, 1.668359281E9, 1.668359329E9, 1.668359377E9, 1.668359425E9, 1.668359473E9, 1.668359521E9, 1.668359569E9, 1.668359617E9, 1.668359665E9, 1.668359713E9, 1.668359761E9, 1.668359809E9, 1.668359857E9, 1.668359905E9, 1.668359953E9, 1.668360001E9, 1.668360049E9, 1.668360097E9, 1.668360145E9, 1.668360193E9, 1.668360241E9, 1.668360289E9, 1.668360337E9, 1.668360385E9, 1.668360433E9, 1.668360481E9, 1.668360529E9, 1.668360577E9, 1.668360625E9, 1.668360673E9, 1.668360721E9, 1.668360769E9, 1.66836108E9, 1.66836126E9, 1.668366939E9, 1.668366987E9, 1.668367035E9, 1.668367083E9, 1.668367131E9, 1.668367179E9, 1.668367227E9, 1.668367275E9, 1.668367323E9, 1.668367371E9, 1.668367419E9, 1.668367467E9, 1.668367515E9, 1.668367563E9, 1.668367611E9, 1.668367659E9, 1.668367707E9, 1.668367755E9, 1.668367803E9, 1.668367851E9, 1.668367899E9, 1.668367947E9, 1.668367995E9, 1.668368043E9, 1.668368091E9, 1.668368139E9, 1.668368187E9, 1.668368235E9, 1.668368283E9, 1.668368331E9, 1.668368379E9, 1.668368427E9, 1.668368475E9, 1.668368523E9, 1.668368571E9, 1.668368619E9, 1.668368667E9, 1.668368715E9, 1.668368763E9, 1.668368811E9, 1.668368859E9, 1.668368907E9, 1.668368955E9, 1.668369003E9, 1.668369051E9, 1.668369099E9, 1.668369147E9, 1.668369195E9, 1.668369243E9, 1.668369291E9, 1.668369339E9, 1.668369387E9, 1.668369435E9, 1.668369483E9, 1.668369531E9, 1.668369579E9, 1.668369627E9, 1.668369675E9, 1.668369723E9, 1.668369771E9, 1.668369819E9, 1.668369867E9, 1.668369915E9, 1.668369963E9, 1.668370011E9, 1.668370059E9, 1.668370107E9, 1.668370155E9, 1.668370203E9, 1.668370251E9, 1.668370299E9, 1.66837068E9, 1.66837086E9, 1.668376572E9, 1.66837662E9, 1.668376668E9, 1.668376716E9, 1.668376764E9, 1.668376812E9, 1.66837686E9, 1.668376908E9, 1.668376956E9, 1.668377004E9, 1.668377052E9, 1.6683771E9, 1.668377148E9, 1.668377196E9, 1.668377244E9, 1.668377292E9, 1.66837734E9, 1.668377388E9, 1.668377436E9, 1.668377484E9, 1.668377532E9, 1.66837758E9, 1.668377628E9, 1.668377676E9, 1.668377724E9, 1.668377772E9, 1.66837782E9, 1.668377868E9, 1.668377916E9, 1.668377964E9, 1.668378012E9, 1.66837806E9, 1.668378108E9, 1.668378156E9, 1.668378204E9, 1.668378252E9, 1.6683783E9, 1.668378348E9, 1.668378396E9, 1.668378444E9, 1.668378492E9, 1.66837854E9, 1.668378588E9, 1.668378636E9, 1.668378684E9, 1.668378732E9, 1.66837878E9, 1.668378828E9, 1.668378876E9, 1.668378924E9, 1.668378972E9, 1.66837902E9, 1.668379068E9, 1.668379116E9, 1.668379164E9, 1.668379212E9, 1.66837926E9, 1.668379308E9, 1.668379356E9, 1.668379404E9, 1.668379452E9, 1.6683795E9, 1.668379548E9, 1.668379596E9, 1.668379644E9, 1.668379692E9, 1.66837974E9, 1.668379788E9, 1.668379836E9, 1.668379884E9, 1.668379932E9, 1.66837998E9, 1.66838028E9, 1.66838046E9, 1.668386198E9, 1.668386246E9, 1.668386294E9, 1.668386342E9, 1.66838639E9, 1.668386438E9, 1.668386486E9, 1.668386534E9, 1.668386582E9, 1.66838663E9, 1.668386678E9, 1.668386726E9, 1.668386774E9, 1.668386822E9, 1.66838687E9, 1.668386918E9, 1.668386966E9, 1.668387014E9, 1.668387062E9, 1.66838711E9, 1.668387158E9, 1.668387206E9, 1.668387254E9, 1.668387302E9, 1.66838735E9, 1.668387398E9, 1.668387446E9, 1.668387494E9, 1.668387542E9, 1.66838759E9, 1.668387638E9, 1.668387686E9, 1.668387734E9, 1.668387782E9, 1.66838783E9, 1.668387878E9, 1.668387926E9, 1.668387974E9, 1.668388022E9, 1.66838807E9, 1.668388118E9, 1.668388166E9, 1.668388214E9, 1.668388262E9, 1.66838831E9, 1.668388358E9, 1.668388406E9, 1.668388454E9, 1.668388502E9, 1.66838855E9, 1.668388598E9, 1.668388646E9, 1.668388694E9, 1.668388742E9, 1.66838879E9, 1.668388838E9, 1.668388886E9, 1.668388934E9, 1.668388982E9, 1.66838903E9, 1.668389078E9, 1.668389126E9, 1.668389174E9, 1.668389222E9, 1.66838927E9, 1.668389318E9, 1.668389366E9, 1.668389414E9, 1.668389462E9, 1.66838951E9, 1.668389558E9, 1.668389606E9, 1.668389654E9, 1.668389702E9, 1.66838975E9, 1.66839E9, 1.66839024E9, 1.668396106E9, 1.668396154E9, 1.668396202E9, 1.66839625E9, 1.668396298E9, 1.668396346E9, 1.668396394E9, 1.668396442E9, 1.66839649E9, 1.668396538E9, 1.668396586E9, 1.668396634E9, 1.668396682E9, 1.66839673E9, 1.668396778E9, 1.668396826E9, 1.668396874E9, 1.668396922E9, 1.66839697E9, 1.668397018E9, 1.668397066E9, 1.668397114E9, 1.668397162E9, 1.66839721E9, 1.668397258E9, 1.668397306E9, 1.668397354E9, 1.668397402E9, 1.66839745E9, 1.668397498E9, 1.668397546E9, 1.668397594E9, 1.668397642E9, 1.66839769E9, 1.668397738E9, 1.668397786E9, 1.668397834E9, 1.668397882E9, 1.66839793E9, 1.668397978E9, 1.668398026E9, 1.668398074E9, 1.668398122E9, 1.66839817E9, 1.668398218E9, 1.668398266E9, 1.668398314E9, 1.668398362E9, 1.66839841E9, 1.668398458E9, 1.668398506E9, 1.668398554E9, 1.668398602E9, 1.66839865E9, 1.668398698E9, 1.668398746E9, 1.668398794E9, 1.668398842E9, 1.66839889E9, 1.668398938E9, 1.668398986E9, 1.668399034E9, 1.668399082E9, 1.66839913E9, 1.668399178E9, 1.668399226E9, 1.668399274E9, 1.668399322E9, 1.66839937E9, 1.66839978E9, 1.66839996E9, 1.668405554E9, 1.668405602E9, 1.66840565E9, 1.668405698E9, 1.668405746E9, 1.668405794E9, 1.668405842E9, 1.66840589E9, 1.668405938E9, 1.668405986E9, 1.668406034E9, 1.668406082E9, 1.66840613E9, 1.668406178E9, 1.668406226E9, 1.668406274E9, 1.668406322E9, 1.66840637E9, 1.668406418E9, 1.668406466E9, 1.668406514E9, 1.668406562E9, 1.66840661E9, 1.668406658E9, 1.668406706E9, 1.668406754E9, 1.668406802E9, 1.66840685E9, 1.668406898E9, 1.668406946E9, 1.668406994E9, 1.668407042E9, 1.66840709E9, 1.668407138E9, 1.668407186E9, 1.668407234E9, 1.668407282E9, 1.66840733E9, 1.668407378E9, 1.668407426E9, 1.668407474E9, 1.668407522E9, 1.66840757E9, 1.668407618E9, 1.668407666E9, 1.668407714E9, 1.668407762E9, 1.66840781E9, 1.668407858E9, 1.668407906E9, 1.668407954E9, 1.668408002E9, 1.66840805E9, 1.668408098E9, 1.668408146E9, 1.668408194E9, 1.668408242E9, 1.66840829E9, 1.668408338E9, 1.668408386E9, 1.668408434E9, 1.668408482E9, 1.66840853E9, 1.668408578E9, 1.668408626E9, 1.668408674E9, 1.668408722E9, 1.66840877E9, 1.66840908E9, 1.66840926E9, 1.668415308E9, 1.668415356E9, 1.668415404E9, 1.668415452E9, 1.6684155E9, 1.668415548E9, 1.668415596E9, 1.668415644E9, 1.668415692E9, 1.66841574E9, 1.668415788E9, 1.668415836E9, 1.668415884E9, 1.668415932E9, 1.66841598E9, 1.668416028E9, 1.668416076E9, 1.668416124E9, 1.668416172E9, 1.66841622E9, 1.668416268E9, 1.668416316E9, 1.668416364E9, 1.668416412E9, 1.66841646E9, 1.668416508E9, 1.668416556E9, 1.668416604E9, 1.668416652E9, 1.6684167E9, 1.668416748E9, 1.668416796E9, 1.668416844E9, 1.668416892E9, 1.66841694E9, 1.668416988E9, 1.668417036E9, 1.668417084E9, 1.668417132E9, 1.66841718E9, 1.668417228E9, 1.668417276E9, 1.668417324E9, 1.668417372E9, 1.66841742E9, 1.668417468E9, 1.668417516E9, 1.668417564E9, 1.668417612E9, 1.66841766E9, 1.668417708E9, 1.668417756E9, 1.668417804E9, 1.668417852E9, 1.6684179E9, 1.668417948E9, 1.668417996E9, 1.668418044E9, 1.668418092E9, 1.66841814E9, 1.668418188E9, 1.668418236E9, 1.668418284E9, 1.668418332E9, 1.66841838E9, 1.668418428E9, 1.668418476E9, 1.668418524E9, 1.668418572E9, 1.66841862E9, 1.66841892E9, 1.6684191E9, 1.668424873E9, 1.668424921E9, 1.668424969E9, 1.668425017E9, 1.668425065E9, 1.668425113E9, 1.668425161E9, 1.668425209E9, 1.668425257E9, 1.668425305E9, 1.668425353E9, 1.668425401E9, 1.668425449E9, 1.668425497E9, 1.668425545E9, 1.668425593E9, 1.668425641E9, 1.668425689E9, 1.668425737E9, 1.668425785E9, 1.668425833E9, 1.668425881E9, 1.668425929E9, 1.668425977E9, 1.668426025E9, 1.668426073E9, 1.668426121E9, 1.668426169E9, 1.668426217E9, 1.668426265E9, 1.668426313E9, 1.668426361E9, 1.668426409E9, 1.668426457E9, 1.668426505E9, 1.668426553E9, 1.668426601E9, 1.668426649E9, 1.668426697E9, 1.668426745E9, 1.668426793E9, 1.668426841E9, 1.668426889E9, 1.668426937E9, 1.668426985E9, 1.668427033E9, 1.668427081E9, 1.668427129E9, 1.668427177E9, 1.668427225E9, 1.668427273E9, 1.668427321E9, 1.668427369E9, 1.668427417E9, 1.668427465E9, 1.668427513E9, 1.668427561E9, 1.668427609E9, 1.668427657E9, 1.668427705E9, 1.668427753E9, 1.668427801E9, 1.668427849E9, 1.668427897E9, 1.668427945E9, 1.668427993E9, 1.668428041E9, 1.668428089E9, 1.6684284E9, 1.66842858E9, 1.668434533E9, 1.668434581E9, 1.668434629E9, 1.668434677E9, 1.668434725E9, 1.668434773E9, 1.668434821E9, 1.668434869E9, 1.668434917E9, 1.668434965E9, 1.668435013E9, 1.668435061E9, 1.668435109E9, 1.668435157E9, 1.668435205E9, 1.668435253E9, 1.668435301E9, 1.668435349E9, 1.668435397E9, 1.668435445E9, 1.668435493E9, 1.668435541E9, 1.668435589E9, 1.668435637E9, 1.668435685E9, 1.668435733E9, 1.668435781E9, 1.668435829E9, 1.668435877E9, 1.668435925E9, 1.668435973E9, 1.668436021E9, 1.668436069E9, 1.668436117E9, 1.668436165E9, 1.668436213E9, 1.668436261E9, 1.668436309E9, 1.668436357E9, 1.668436405E9, 1.668436453E9, 1.668436501E9, 1.668436549E9, 1.668436597E9, 1.668436645E9, 1.668436693E9, 1.668436741E9, 1.668436789E9, 1.668436837E9, 1.668436885E9, 1.668436933E9, 1.668436981E9, 1.668437029E9, 1.668437077E9, 1.668437125E9, 1.668437173E9, 1.668437221E9, 1.668437269E9, 1.668437317E9, 1.668437365E9, 1.668437413E9, 1.668437461E9, 1.668437509E9, 1.668437557E9, 1.668437605E9, 1.668437653E9, 1.668437701E9, 1.668437749E9, 1.66843806E9, 1.66843824E9, 1.66844415E9, 1.668444198E9, 1.668444246E9, 1.668444294E9, 1.668444342E9, 1.66844439E9, 1.668444438E9, 1.668444486E9, 1.668444534E9, 1.668444582E9, 1.66844463E9, 1.668444678E9, 1.668444726E9, 1.668444774E9, 1.668444822E9, 1.66844487E9, 1.668444918E9, 1.668444966E9, 1.668445014E9, 1.668445062E9, 1.66844511E9, 1.668445158E9, 1.668445206E9, 1.668445254E9, 1.668445302E9, 1.66844535E9, 1.668445398E9, 1.668445446E9, 1.668445494E9, 1.668445542E9, 1.66844559E9, 1.668445638E9, 1.668445686E9, 1.668445734E9, 1.668445782E9, 1.66844583E9, 1.668445878E9, 1.668445926E9, 1.668445974E9, 1.668446022E9, 1.66844607E9, 1.668446118E9, 1.668446166E9, 1.668446214E9, 1.668446262E9, 1.66844631E9, 1.668446358E9, 1.668446406E9, 1.668446454E9, 1.668446502E9, 1.66844655E9, 1.668446598E9, 1.668446646E9, 1.668446694E9, 1.668446742E9, 1.66844679E9, 1.668446838E9, 1.668446886E9, 1.668446934E9, 1.668446982E9, 1.66844703E9, 1.668447078E9, 1.668447126E9, 1.668447174E9, 1.668447222E9, 1.66844727E9, 1.668447318E9, 1.668447366E9, 1.668447414E9, 1.668447462E9, 1.66844751E9, 1.66844778E9, 1.66844796E9, 1.668453821E9, 1.668453869E9, 1.668453917E9, 1.668453965E9, 1.668454013E9, 1.668454061E9, 1.668454109E9, 1.668454157E9, 1.668454205E9, 1.668454253E9, 1.668454301E9, 1.668454349E9, 1.668454397E9, 1.668454445E9, 1.668454493E9, 1.668454541E9, 1.668454589E9, 1.668454637E9, 1.668454685E9, 1.668454733E9, 1.668454781E9, 1.668454829E9, 1.668454877E9, 1.668454925E9, 1.668454973E9, 1.668455021E9, 1.668455069E9, 1.668455117E9, 1.668455165E9, 1.668455213E9, 1.668455261E9, 1.668455309E9, 1.668455357E9, 1.668455405E9, 1.668455453E9, 1.668455501E9, 1.668455549E9, 1.668455597E9, 1.668455645E9, 1.668455693E9, 1.668455741E9, 1.668455789E9, 1.668455837E9, 1.668455885E9, 1.668455933E9, 1.668455981E9, 1.668456029E9, 1.668456077E9, 1.668456125E9, 1.668456173E9, 1.668456221E9, 1.668456269E9, 1.668456317E9, 1.668456365E9, 1.668456413E9, 1.668456461E9, 1.668456509E9, 1.668456557E9, 1.668456605E9, 1.668456653E9, 1.668456701E9, 1.668456749E9, 1.668456797E9, 1.668456845E9, 1.668456893E9, 1.668456941E9, 1.668456989E9, 1.66845732E9, 1.6684575E9, 1.668463243E9, 1.668463291E9, 1.668463339E9, 1.668463387E9, 1.668463435E9, 1.668463483E9, 1.668463531E9, 1.668463579E9, 1.668463627E9, 1.668463675E9, 1.668463723E9, 1.668463771E9, 1.668463819E9, 1.668463867E9, 1.668463915E9, 1.668463963E9, 1.668464011E9, 1.668464059E9, 1.668464107E9, 1.668464155E9, 1.668464203E9, 1.668464251E9, 1.668464299E9, 1.668464347E9, 1.668464395E9, 1.668464443E9, 1.668464491E9, 1.668464539E9, 1.668464587E9, 1.668464635E9, 1.668464683E9, 1.668464731E9, 1.668464779E9, 1.668464827E9, 1.668464875E9, 1.668464923E9, 1.668464971E9, 1.668465019E9, 1.668465067E9, 1.668465115E9, 1.668465163E9, 1.668465211E9, 1.668465259E9, 1.668465307E9, 1.668465355E9, 1.668465403E9, 1.668465451E9, 1.668465499E9, 1.668465547E9, 1.668465595E9, 1.668465643E9, 1.668465691E9, 1.668465739E9, 1.668465787E9, 1.668465835E9, 1.668465883E9, 1.668465931E9, 1.668465979E9, 1.668466027E9, 1.668466075E9, 1.668466123E9, 1.668466171E9, 1.668466219E9, 1.668466267E9, 1.668466315E9, 1.668466363E9, 1.668466411E9, 1.668466459E9, 1.66846674E9, 1.66846692E9, 1.668472615E9, 1.668472663E9, 1.668472711E9, 1.668472759E9, 1.668472807E9, 1.668472855E9, 1.668472903E9, 1.668472951E9, 1.668472999E9, 1.668473047E9, 1.668473095E9, 1.668473143E9, 1.668473191E9, 1.668473239E9, 1.668473287E9, 1.668473335E9, 1.668473383E9, 1.668473431E9, 1.668473479E9, 1.668473527E9, 1.668473575E9, 1.668473623E9, 1.668473671E9, 1.668473719E9, 1.668473767E9, 1.668473815E9, 1.668473863E9, 1.668473911E9, 1.668473959E9, 1.668474007E9, 1.668474055E9, 1.668474103E9, 1.668474151E9, 1.668474199E9, 1.668474247E9, 1.668474295E9, 1.668474343E9, 1.668474391E9, 1.668474439E9, 1.668474487E9, 1.668474535E9, 1.668474583E9, 1.668474631E9, 1.668474679E9, 1.668474727E9, 1.668474775E9, 1.668474823E9, 1.668474871E9, 1.668474919E9, 1.668474967E9, 1.668475015E9, 1.668475063E9, 1.668475111E9, 1.668475159E9, 1.668475207E9, 1.668475255E9, 1.668475303E9, 1.668475351E9, 1.668475399E9, 1.668475447E9, 1.668475495E9, 1.668475543E9, 1.668475591E9, 1.668475639E9, 1.668475687E9, 1.668475735E9, 1.668475783E9, 1.668475831E9, 1.668475879E9, 1.66847616E9, 1.66847634E9, 1.668481976E9, 1.668482024E9, 1.668482072E9, 1.66848212E9, 1.668482168E9, 1.668482216E9, 1.668482264E9, 1.668482312E9, 1.66848236E9, 1.668482408E9, 1.668482456E9, 1.668482504E9, 1.668482552E9, 1.6684826E9, 1.668482648E9, 1.668482696E9, 1.668482744E9, 1.668482792E9, 1.66848284E9, 1.668482888E9, 1.668482936E9, 1.668482984E9, 1.668483032E9, 1.66848308E9, 1.668483128E9, 1.668483176E9, 1.668483224E9, 1.668483272E9, 1.66848332E9, 1.668483368E9, 1.668483416E9, 1.668483464E9, 1.668483512E9, 1.66848356E9, 1.668483608E9, 1.668483656E9, 1.668483704E9, 1.668483752E9, 1.6684838E9, 1.668483848E9, 1.668483896E9, 1.668483944E9, 1.668483992E9, 1.66848404E9, 1.668484088E9, 1.668484136E9, 1.668484184E9, 1.668484232E9, 1.66848428E9, 1.668484328E9, 1.668484376E9, 1.668484424E9, 1.668484472E9, 1.66848452E9, 1.668484568E9, 1.668484616E9, 1.668484664E9, 1.668484712E9, 1.66848476E9, 1.668484808E9, 1.668484856E9, 1.668484904E9, 1.668484952E9, 1.668485E9, 1.668485048E9, 1.668485096E9, 1.668485144E9, 1.668485192E9, 1.66848524E9, 1.66848558E9, 1.66848576E9, 1.668491391E9, 1.668491439E9, 1.668491487E9, 1.668491535E9, 1.668491583E9, 1.668491631E9, 1.668491679E9, 1.668491727E9, 1.668491775E9, 1.668491823E9, 1.668491871E9, 1.668491919E9, 1.668491967E9, 1.668492015E9, 1.668492063E9, 1.668492111E9, 1.668492159E9, 1.668492207E9, 1.668492255E9, 1.668492303E9, 1.668492351E9, 1.668492399E9, 1.668492447E9, 1.668492495E9, 1.668492543E9, 1.668492591E9, 1.668492639E9, 1.668492687E9, 1.668492735E9, 1.668492783E9, 1.668492831E9, 1.668492879E9, 1.668492927E9, 1.668492975E9, 1.668493023E9, 1.668493071E9, 1.668493119E9, 1.668493167E9, 1.668493215E9, 1.668493263E9, 1.668493311E9, 1.668493359E9, 1.668493407E9, 1.668493455E9, 1.668493503E9, 1.668493551E9, 1.668493599E9, 1.668493647E9, 1.668493695E9, 1.668493743E9, 1.668493791E9, 1.668493839E9, 1.668493887E9, 1.668493935E9, 1.668493983E9, 1.668494031E9, 1.668494079E9, 1.668494127E9, 1.668494175E9, 1.668494223E9, 1.668494271E9, 1.668494319E9, 1.668494367E9, 1.668494415E9, 1.668494463E9, 1.668494511E9, 1.668494559E9, 1.668494607E9, 1.668494655E9, 1.668494703E9, 1.668494751E9, 1.668494799E9, 1.66849506E9, 1.66849524E9, 1.668500926E9, 1.668500974E9, 1.668501022E9, 1.66850107E9, 1.668501118E9, 1.668501166E9, 1.668501214E9, 1.668501262E9, 1.66850131E9, 1.668501358E9, 1.668501406E9, 1.668501454E9, 1.668501502E9, 1.66850155E9, 1.668501598E9, 1.668501646E9, 1.668501694E9, 1.668501742E9, 1.66850179E9, 1.668501838E9, 1.668501886E9, 1.668501934E9, 1.668501982E9, 1.66850203E9, 1.668502078E9, 1.668502126E9, 1.668502174E9, 1.668502222E9, 1.66850227E9, 1.668502318E9, 1.668502366E9, 1.668502414E9, 1.668502462E9, 1.66850251E9, 1.668502558E9, 1.668502606E9, 1.668502654E9, 1.668502702E9, 1.66850275E9, 1.668502798E9, 1.668502846E9, 1.668502894E9, 1.668502942E9, 1.66850299E9, 1.668503038E9, 1.668503086E9, 1.668503134E9, 1.668503182E9, 1.66850323E9, 1.668503278E9, 1.668503326E9, 1.668503374E9, 1.668503422E9, 1.66850347E9, 1.668503518E9, 1.668503566E9, 1.668503614E9, 1.668503662E9, 1.66850371E9, 1.668503758E9, 1.668503806E9, 1.668503854E9, 1.668503902E9, 1.66850395E9, 1.668503998E9, 1.668504046E9, 1.668504094E9, 1.668504142E9, 1.66850419E9, 1.66850448E9, 1.66850466E9, 1.668510401E9, 1.668510449E9, 1.668510497E9, 1.668510545E9, 1.668510593E9, 1.668510641E9, 1.668510689E9, 1.668510737E9, 1.668510785E9, 1.668510833E9, 1.668510881E9, 1.668510929E9, 1.668510977E9, 1.668511025E9, 1.668511073E9, 1.668511121E9, 1.668511169E9, 1.668511217E9, 1.668511265E9, 1.668511313E9, 1.668511361E9, 1.668511409E9, 1.668511457E9, 1.668511505E9, 1.668511553E9, 1.668511601E9, 1.668511649E9, 1.668511697E9, 1.668511745E9, 1.668511793E9, 1.668511841E9, 1.668511889E9, 1.668511937E9, 1.668511985E9, 1.668512033E9, 1.668512081E9, 1.668512129E9, 1.668512177E9, 1.668512225E9, 1.668512273E9, 1.668512321E9, 1.668512369E9, 1.668512417E9, 1.668512465E9, 1.668512513E9, 1.668512561E9, 1.668512609E9, 1.668512657E9, 1.668512705E9, 1.668512753E9, 1.668512801E9, 1.668512849E9, 1.668512897E9, 1.668512945E9, 1.668512993E9, 1.668513041E9, 1.668513089E9, 1.668513137E9, 1.668513185E9, 1.668513233E9, 1.668513281E9, 1.668513329E9, 1.668513377E9, 1.668513425E9, 1.668513473E9, 1.668513521E9, 1.668513569E9, 1.668513617E9, 1.668513665E9, 1.668513713E9, 1.668513761E9, 1.668513809E9, 1.66851414E9, 1.66851432E9, 1.668519946E9, 1.668519994E9, 1.668520042E9, 1.66852009E9, 1.668520138E9, 1.668520186E9, 1.668520234E9, 1.668520282E9, 1.66852033E9, 1.668520378E9, 1.668520426E9, 1.668520474E9, 1.668520522E9, 1.66852057E9, 1.668520618E9, 1.668520666E9, 1.668520714E9, 1.668520762E9, 1.66852081E9, 1.668520858E9, 1.668520906E9, 1.668520954E9, 1.668521002E9, 1.66852105E9, 1.668521098E9, 1.668521146E9, 1.668521194E9, 1.668521242E9, 1.66852129E9, 1.668521338E9, 1.668521386E9, 1.668521434E9, 1.668521482E9, 1.66852153E9, 1.668521578E9, 1.668521626E9, 1.668521674E9, 1.668521722E9, 1.66852177E9, 1.668521818E9, 1.668521866E9, 1.668521914E9, 1.668521962E9, 1.66852201E9, 1.668522058E9, 1.668522106E9, 1.668522154E9, 1.668522202E9, 1.66852225E9, 1.668522298E9, 1.668522346E9, 1.668522394E9, 1.668522442E9, 1.66852249E9, 1.668522538E9, 1.668522586E9, 1.668522634E9, 1.668522682E9, 1.66852273E9, 1.668522778E9, 1.668522826E9, 1.668522874E9, 1.668522922E9, 1.66852297E9, 1.668523018E9, 1.668523066E9, 1.668523114E9, 1.668523162E9, 1.66852321E9, 1.6685235E9, 1.66852368E9, 1.668529713E9, 1.668529761E9, 1.668529809E9, 1.668529857E9, 1.668529905E9, 1.668529953E9, 1.668530001E9, 1.668530049E9, 1.668530097E9, 1.668530145E9, 1.668530193E9, 1.668530241E9, 1.668530289E9, 1.668530337E9, 1.668530385E9, 1.668530433E9, 1.668530481E9, 1.668530529E9, 1.668530577E9, 1.668530625E9, 1.668530673E9, 1.668530721E9, 1.668530769E9, 1.668530817E9, 1.668530865E9, 1.668530913E9, 1.668530961E9, 1.668531009E9, 1.668531057E9, 1.668531105E9, 1.668531153E9, 1.668531201E9, 1.668531249E9, 1.668531297E9, 1.668531345E9, 1.668531393E9, 1.668531441E9, 1.668531489E9, 1.668531537E9, 1.668531585E9, 1.668531633E9, 1.668531681E9, 1.668531729E9, 1.668531777E9, 1.668531825E9, 1.668531873E9, 1.668531921E9, 1.668531969E9, 1.668532017E9, 1.668532065E9, 1.668532113E9, 1.668532161E9, 1.668532209E9, 1.668532257E9, 1.668532305E9, 1.668532353E9, 1.668532401E9, 1.668532449E9, 1.668532497E9, 1.668532545E9, 1.668532593E9, 1.668532641E9, 1.668532689E9, 1.668532737E9, 1.668532785E9, 1.668532833E9, 1.668532881E9, 1.668532929E9, 1.66853322E9, 1.6685334E9, 1.668539355E9, 1.668539403E9, 1.668539451E9, 1.668539499E9, 1.668539547E9, 1.668539595E9, 1.668539643E9, 1.668539691E9, 1.668539739E9, 1.668539787E9, 1.668539835E9, 1.668539883E9, 1.668539931E9, 1.668539979E9, 1.668540027E9, 1.668540075E9, 1.668540123E9, 1.668540171E9, 1.668540219E9, 1.668540267E9, 1.668540315E9, 1.668540363E9, 1.668540411E9, 1.668540459E9, 1.668540507E9, 1.668540555E9, 1.668540603E9, 1.668540651E9, 1.668540699E9, 1.668540747E9, 1.668540795E9, 1.668540843E9, 1.668540891E9, 1.668540939E9, 1.668540987E9, 1.668541035E9, 1.668541083E9, 1.668541131E9, 1.668541179E9, 1.668541227E9, 1.668541275E9, 1.668541323E9, 1.668541371E9, 1.668541419E9, 1.668541467E9, 1.668541515E9, 1.668541563E9, 1.668541611E9, 1.668541659E9, 1.668541707E9, 1.668541755E9, 1.668541803E9, 1.668541851E9, 1.668541899E9, 1.668541947E9, 1.668541995E9, 1.668542043E9, 1.668542091E9, 1.668542139E9, 1.668542187E9, 1.668542235E9, 1.668542283E9, 1.668542331E9, 1.668542379E9, 1.668542427E9, 1.668542475E9, 1.668542523E9, 1.668542571E9, 1.668542619E9, 1.668543E9, 1.66854318E9, 1.668548855E9, 1.668548903E9, 1.668548951E9, 1.668548999E9, 1.668549047E9, 1.668549095E9, 1.668549143E9, 1.668549191E9, 1.668549239E9, 1.668549287E9, 1.668549335E9, 1.668549383E9, 1.668549431E9, 1.668549479E9, 1.668549527E9, 1.668549575E9, 1.668549623E9, 1.668549671E9, 1.668549719E9, 1.668549767E9, 1.668549815E9, 1.668549863E9, 1.668549911E9, 1.668549959E9, 1.668550007E9, 1.668550055E9, 1.668550103E9, 1.668550151E9, 1.668550199E9, 1.668550247E9, 1.668550295E9, 1.668550343E9, 1.668550391E9, 1.668550439E9, 1.668550487E9, 1.668550535E9, 1.668550583E9, 1.668550631E9, 1.668550679E9, 1.668550727E9, 1.668550775E9, 1.668550823E9, 1.668550871E9, 1.668550919E9, 1.668550967E9, 1.668551015E9, 1.668551063E9, 1.668551111E9, 1.668551159E9, 1.668551207E9, 1.668551255E9, 1.668551303E9, 1.668551351E9, 1.668551399E9, 1.668551447E9, 1.668551495E9, 1.668551543E9, 1.668551591E9, 1.668551639E9, 1.668551687E9, 1.668551735E9, 1.668551783E9, 1.668551831E9, 1.668551879E9, 1.668551927E9, 1.668551975E9, 1.668552023E9, 1.668552071E9, 1.668552119E9, 1.66855242E9, 1.6685526E9, 1.668558444E9, 1.668558492E9, 1.66855854E9, 1.668558588E9, 1.668558636E9, 1.668558684E9, 1.668558732E9, 1.66855878E9, 1.668558828E9, 1.668558876E9, 1.668558924E9, 1.668558972E9, 1.66855902E9, 1.668559068E9, 1.668559116E9, 1.668559164E9, 1.668559212E9, 1.66855926E9, 1.668559308E9, 1.668559356E9, 1.668559404E9, 1.668559452E9, 1.6685595E9, 1.668559548E9, 1.668559596E9, 1.668559644E9, 1.668559692E9, 1.66855974E9, 1.668559788E9, 1.668559836E9, 1.668559884E9, 1.668559932E9, 1.66855998E9, 1.668560028E9, 1.668560076E9, 1.668560124E9, 1.668560172E9, 1.66856022E9, 1.668560268E9, 1.668560316E9, 1.668560364E9, 1.668560412E9, 1.66856046E9, 1.668560508E9, 1.668560556E9, 1.668560604E9, 1.668560652E9, 1.6685607E9, 1.668560748E9, 1.668560796E9, 1.668560844E9, 1.668560892E9, 1.66856094E9, 1.668560988E9, 1.668561036E9, 1.668561084E9, 1.668561132E9, 1.66856118E9, 1.668561228E9, 1.668561276E9, 1.668561324E9, 1.668561372E9, 1.66856142E9, 1.668561468E9, 1.668561516E9, 1.668561564E9, 1.668561612E9, 1.66856166E9, 1.66856196E9, 1.66856214E9, 1.668567836E9, 1.668567884E9, 1.668567932E9, 1.66856798E9, 1.668568028E9, 1.668568076E9, 1.668568124E9, 1.668568172E9, 1.66856822E9, 1.668568268E9, 1.668568316E9, 1.668568364E9, 1.668568412E9, 1.66856846E9, 1.668568508E9, 1.668568556E9, 1.668568604E9, 1.668568652E9, 1.6685687E9, 1.668568748E9, 1.668568796E9, 1.668568844E9, 1.668568892E9, 1.66856894E9, 1.668568988E9, 1.668569036E9, 1.668569084E9, 1.668569132E9, 1.66856918E9, 1.668569228E9, 1.668569276E9, 1.668569324E9, 1.668569372E9, 1.66856942E9, 1.668569468E9, 1.668569516E9, 1.668569564E9, 1.668569612E9, 1.66856966E9, 1.668569708E9, 1.668569756E9, 1.668569804E9, 1.668569852E9, 1.6685699E9, 1.668569948E9, 1.668569996E9, 1.668570044E9, 1.668570092E9, 1.66857014E9, 1.668570188E9, 1.668570236E9, 1.668570284E9, 1.668570332E9, 1.66857038E9, 1.668570428E9, 1.668570476E9, 1.668570524E9, 1.668570572E9, 1.66857062E9, 1.668570668E9, 1.668570716E9, 1.668570764E9, 1.668570812E9, 1.66857086E9, 1.668570908E9, 1.668570956E9, 1.668571004E9, 1.668571052E9, 1.6685711E9, 1.66857144E9, 1.66857162E9, 1.668577359E9, 1.668577407E9, 1.668577455E9, 1.668577503E9, 1.668577551E9, 1.668577599E9, 1.668577647E9, 1.668577695E9, 1.668577743E9, 1.668577791E9, 1.668577839E9, 1.668577887E9, 1.668577935E9, 1.668577983E9, 1.668578031E9, 1.668578079E9, 1.668578127E9, 1.668578175E9, 1.668578223E9, 1.668578271E9, 1.668578319E9, 1.668578367E9, 1.668578415E9, 1.668578463E9, 1.668578511E9, 1.668578559E9, 1.668578607E9, 1.668578655E9, 1.668578703E9, 1.668578751E9, 1.668578799E9, 1.668578847E9, 1.668578895E9, 1.668578943E9, 1.668578991E9, 1.668579039E9, 1.668579087E9, 1.668579135E9, 1.668579183E9, 1.668579231E9, 1.668579279E9, 1.668579327E9, 1.668579375E9, 1.668579423E9, 1.668579471E9, 1.668579519E9, 1.668579567E9, 1.668579615E9, 1.668579663E9, 1.668579711E9, 1.668579759E9, 1.668579807E9, 1.668579855E9, 1.668579903E9, 1.668579951E9, 1.668579999E9, 1.668580047E9, 1.668580095E9, 1.668580143E9, 1.668580191E9, 1.668580239E9, 1.668580287E9, 1.668580335E9, 1.668580383E9, 1.668580431E9, 1.668580479E9, 1.6685808E9, 1.66858098E9, 1.668586829E9, 1.668586877E9, 1.668586925E9, 1.668586973E9, 1.668587021E9, 1.668587069E9, 1.668587117E9, 1.668587165E9, 1.668587213E9, 1.668587261E9, 1.668587309E9, 1.668587357E9, 1.668587405E9, 1.668587453E9, 1.668587501E9, 1.668587549E9, 1.668587597E9, 1.668587645E9, 1.668587693E9, 1.668587741E9, 1.668587789E9, 1.668587837E9, 1.668587885E9, 1.668587933E9, 1.668587981E9, 1.668588029E9, 1.668588077E9, 1.668588125E9, 1.668588173E9, 1.668588221E9, 1.668588269E9, 1.668588317E9, 1.668588365E9, 1.668588413E9, 1.668588461E9, 1.668588509E9, 1.668588557E9, 1.668588605E9, 1.668588653E9, 1.668588701E9, 1.668588749E9, 1.668588797E9, 1.668588845E9, 1.668588893E9, 1.668588941E9, 1.668588989E9, 1.668589037E9, 1.668589085E9, 1.668589133E9, 1.668589181E9, 1.668589229E9, 1.668589277E9, 1.668589325E9, 1.668589373E9, 1.668589421E9, 1.668589469E9, 1.668589517E9, 1.668589565E9, 1.668589613E9, 1.668589661E9, 1.668589709E9, 1.668589757E9, 1.668589805E9, 1.668589853E9, 1.668589901E9, 1.668589949E9, 1.668589997E9, 1.668590045E9, 1.668590093E9, 1.668590141E9, 1.668590189E9, 1.66859058E9, 1.66859076E9, 1.668596358E9, 1.668596406E9, 1.668596454E9, 1.668596502E9, 1.66859655E9, 1.668596598E9, 1.668596646E9, 1.668596694E9, 1.668596742E9, 1.66859679E9, 1.668596838E9, 1.668596886E9, 1.668596934E9, 1.668596982E9, 1.66859703E9, 1.668597078E9, 1.668597126E9, 1.668597174E9, 1.668597222E9, 1.66859727E9, 1.668597318E9, 1.668597366E9, 1.668597414E9, 1.668597462E9, 1.66859751E9, 1.668597558E9, 1.668597606E9, 1.668597654E9, 1.668597702E9, 1.66859775E9, 1.668597798E9, 1.668597846E9, 1.668597894E9, 1.668597942E9, 1.66859799E9, 1.668598038E9, 1.668598086E9, 1.668598134E9, 1.668598182E9, 1.66859823E9, 1.668598278E9, 1.668598326E9, 1.668598374E9, 1.668598422E9, 1.66859847E9, 1.668598518E9, 1.668598566E9, 1.668598614E9, 1.668598662E9, 1.66859871E9, 1.668598758E9, 1.668598806E9, 1.668598854E9, 1.668598902E9, 1.66859895E9, 1.668598998E9, 1.668599046E9, 1.668599094E9, 1.668599142E9, 1.66859919E9, 1.668599238E9, 1.668599286E9, 1.668599334E9, 1.668599382E9, 1.66859943E9, 1.668599478E9, 1.668599526E9, 1.668599574E9, 1.668599622E9, 1.66859967E9, 1.6686E9, 1.66860018E9, 1.668605895E9, 1.668605943E9, 1.668605991E9, 1.668606039E9, 1.668606087E9, 1.668606135E9, 1.668606183E9, 1.668606231E9, 1.668606279E9, 1.668606327E9, 1.668606375E9, 1.668606423E9, 1.668606471E9, 1.668606519E9, 1.668606567E9, 1.668606615E9, 1.668606663E9, 1.668606711E9, 1.668606759E9, 1.668606807E9, 1.668606855E9, 1.668606903E9, 1.668606951E9, 1.668606999E9, 1.668607047E9, 1.668607095E9, 1.668607143E9, 1.668607191E9, 1.668607239E9, 1.668607287E9, 1.668607335E9, 1.668607383E9, 1.668607431E9, 1.668607479E9, 1.668607527E9, 1.668607575E9, 1.668607623E9, 1.668607671E9, 1.668607719E9, 1.668607767E9, 1.668607815E9, 1.668607863E9, 1.668607911E9, 1.668607959E9, 1.668608007E9, 1.668608055E9, 1.668608103E9, 1.668608151E9, 1.668608199E9, 1.668608247E9, 1.668608295E9, 1.668608343E9, 1.668608391E9, 1.668608439E9, 1.668608487E9, 1.668608535E9, 1.668608583E9, 1.668608631E9, 1.668608679E9, 1.668608727E9, 1.668608775E9, 1.668608823E9, 1.668608871E9, 1.668608919E9, 1.668608967E9, 1.668609015E9, 1.668609063E9, 1.668609111E9, 1.668609159E9, 1.66860948E9, 1.66860966E9, 1.668615405E9, 1.668615453E9, 1.668615501E9, 1.668615549E9, 1.668615597E9, 1.668615645E9, 1.668615693E9, 1.668615741E9, 1.668615789E9, 1.668615837E9, 1.668615885E9, 1.668615933E9, 1.668615981E9, 1.668616029E9, 1.668616077E9, 1.668616125E9, 1.668616173E9, 1.668616221E9, 1.668616269E9, 1.668616317E9, 1.668616365E9, 1.668616413E9, 1.668616461E9, 1.668616509E9, 1.668616557E9, 1.668616605E9, 1.668616653E9, 1.668616701E9, 1.668616749E9, 1.668616797E9, 1.668616845E9, 1.668616893E9, 1.668616941E9, 1.668616989E9, 1.668617037E9, 1.668617085E9, 1.668617133E9, 1.668617181E9, 1.668617229E9, 1.668617277E9, 1.668617325E9, 1.668617373E9, 1.668617421E9, 1.668617469E9, 1.668617517E9, 1.668617565E9, 1.668617613E9, 1.668617661E9, 1.668617709E9, 1.668617757E9, 1.668617805E9, 1.668617853E9, 1.668617901E9, 1.668617949E9, 1.668617997E9, 1.668618045E9, 1.668618093E9, 1.668618141E9, 1.668618189E9, 1.668618237E9, 1.668618285E9, 1.668618333E9, 1.668618381E9, 1.668618429E9, 1.668618477E9, 1.668618525E9, 1.668618573E9, 1.668618621E9, 1.668618669E9, 1.66861896E9, 1.66861914E9, 1.668624876E9, 1.668624924E9, 1.668624972E9, 1.66862502E9, 1.668625068E9, 1.668625116E9, 1.668625164E9, 1.668625212E9, 1.66862526E9, 1.668625308E9, 1.668625356E9, 1.668625404E9, 1.668625452E9, 1.6686255E9, 1.668625548E9, 1.668625596E9, 1.668625644E9, 1.668625692E9, 1.66862574E9, 1.668625788E9, 1.668625836E9, 1.668625884E9, 1.668625932E9, 1.66862598E9, 1.668626028E9, 1.668626076E9, 1.668626124E9, 1.668626172E9, 1.66862622E9, 1.668626268E9, 1.668626316E9, 1.668626364E9, 1.668626412E9, 1.66862646E9, 1.668626508E9, 1.668626556E9, 1.668626604E9, 1.668626652E9, 1.6686267E9, 1.668626748E9, 1.668626796E9, 1.668626844E9, 1.668626892E9, 1.66862694E9, 1.668626988E9, 1.668627036E9, 1.668627084E9, 1.668627132E9, 1.66862718E9, 1.668627228E9, 1.668627276E9, 1.668627324E9, 1.668627372E9, 1.66862742E9, 1.668627468E9, 1.668627516E9, 1.668627564E9, 1.668627612E9, 1.66862766E9, 1.668627708E9, 1.668627756E9, 1.668627804E9, 1.668627852E9, 1.6686279E9, 1.668627948E9, 1.668627996E9, 1.668628044E9, 1.668628092E9, 1.66862814E9, 1.668628188E9, 1.668628236E9, 1.668628284E9, 1.668628332E9, 1.66862838E9, 1.66862868E9, 1.66862886E9, 1.66863487E9, 1.668634918E9, 1.668634966E9, 1.668635014E9, 1.668635062E9, 1.66863511E9, 1.668635158E9, 1.668635206E9, 1.668635254E9, 1.668635302E9, 1.66863535E9, 1.668635398E9, 1.668635446E9, 1.668635494E9, 1.668635542E9, 1.66863559E9, 1.668635638E9, 1.668635686E9, 1.668635734E9, 1.668635782E9, 1.66863583E9, 1.668635878E9, 1.668635926E9, 1.668635974E9, 1.668636022E9, 1.66863607E9, 1.668636118E9, 1.668636166E9, 1.668636214E9, 1.668636262E9, 1.66863631E9, 1.668636358E9, 1.668636406E9, 1.668636454E9, 1.668636502E9, 1.66863655E9, 1.668636598E9, 1.668636646E9, 1.668636694E9, 1.668636742E9, 1.66863679E9, 1.668636838E9, 1.668636886E9, 1.668636934E9, 1.668636982E9, 1.66863703E9, 1.668637078E9, 1.668637126E9, 1.668637174E9, 1.668637222E9, 1.66863727E9, 1.668637318E9, 1.668637366E9, 1.668637414E9, 1.668637462E9, 1.66863751E9, 1.668637558E9, 1.668637606E9, 1.668637654E9, 1.668637702E9, 1.66863775E9, 1.668637798E9, 1.668637846E9, 1.668637894E9, 1.668637942E9, 1.66863799E9, 1.668638038E9, 1.668638086E9, 1.668638134E9, 1.668638182E9, 1.66863823E9, 1.66863858E9, 1.66863876E9, 1.668644572E9, 1.66864462E9, 1.668644668E9, 1.668644716E9, 1.668644764E9, 1.668644812E9, 1.66864486E9, 1.668644908E9, 1.668644956E9, 1.668645004E9, 1.668645052E9, 1.6686451E9, 1.668645148E9, 1.668645196E9, 1.668645244E9, 1.668645292E9, 1.66864534E9, 1.668645388E9, 1.668645436E9, 1.668645484E9, 1.668645532E9, 1.66864558E9, 1.668645628E9, 1.668645676E9, 1.668645724E9, 1.668645772E9, 1.66864582E9, 1.668645868E9, 1.668645916E9, 1.668645964E9, 1.668646012E9, 1.66864606E9, 1.668646108E9, 1.668646156E9, 1.668646204E9, 1.668646252E9, 1.6686463E9, 1.668646348E9, 1.668646396E9, 1.668646444E9, 1.668646492E9, 1.66864654E9, 1.668646588E9, 1.668646636E9, 1.668646684E9, 1.668646732E9, 1.66864678E9, 1.668646828E9, 1.668646876E9, 1.668646924E9, 1.668646972E9, 1.66864702E9, 1.668647068E9, 1.668647116E9, 1.668647164E9, 1.668647212E9, 1.66864726E9, 1.668647308E9, 1.668647356E9, 1.668647404E9, 1.668647452E9, 1.6686475E9, 1.668647548E9, 1.668647596E9, 1.668647644E9, 1.668647692E9, 1.66864774E9, 1.668647788E9, 1.668647836E9, 1.668647884E9, 1.668647932E9, 1.66864798E9, 1.66864824E9, 1.66864848E9, 1.668654302E9, 1.66865435E9, 1.668654398E9, 1.668654446E9, 1.668654494E9, 1.668654542E9, 1.66865459E9, 1.668654638E9, 1.668654686E9, 1.668654734E9, 1.668654782E9, 1.66865483E9, 1.668654878E9, 1.668654926E9, 1.668654974E9, 1.668655022E9, 1.66865507E9, 1.668655118E9, 1.668655166E9, 1.668655214E9, 1.668655262E9, 1.66865531E9, 1.668655358E9, 1.668655406E9, 1.668655454E9, 1.668655502E9, 1.66865555E9, 1.668655598E9, 1.668655646E9, 1.668655694E9, 1.668655742E9, 1.66865579E9, 1.668655838E9, 1.668655886E9, 1.668655934E9, 1.668655982E9, 1.66865603E9, 1.668656078E9, 1.668656126E9, 1.668656174E9, 1.668656222E9, 1.66865627E9, 1.668656318E9, 1.668656366E9, 1.668656414E9, 1.668656462E9, 1.66865651E9, 1.668656558E9, 1.668656606E9, 1.668656654E9, 1.668656702E9, 1.66865675E9, 1.668656798E9, 1.668656846E9, 1.668656894E9, 1.668656942E9, 1.66865699E9, 1.668657038E9, 1.668657086E9, 1.668657134E9, 1.668657182E9, 1.66865723E9, 1.668657278E9, 1.668657326E9, 1.668657374E9, 1.668657422E9, 1.66865747E9, 1.668657518E9, 1.668657566E9, 1.668657614E9, 1.668657662E9, 1.66865771E9, 1.668657758E9, 1.668657806E9, 1.668657854E9, 1.668657902E9, 1.66865795E9, 1.66865832E9, 1.6686585E9, 1.668664287E9, 1.668664335E9, 1.668664383E9, 1.668664431E9, 1.668664479E9, 1.668664527E9, 1.668664575E9, 1.668664623E9, 1.668664671E9, 1.668664719E9, 1.668664767E9, 1.668664815E9, 1.668664863E9, 1.668664911E9, 1.668664959E9, 1.668665007E9, 1.668665055E9, 1.668665103E9, 1.668665151E9, 1.668665199E9, 1.668665247E9, 1.668665295E9, 1.668665343E9, 1.668665391E9, 1.668665439E9, 1.668665487E9, 1.668665535E9, 1.668665583E9, 1.668665631E9, 1.668665679E9, 1.668665727E9, 1.668665775E9, 1.668665823E9, 1.668665871E9, 1.668665919E9, 1.668665967E9, 1.668666015E9, 1.668666063E9, 1.668666111E9, 1.668666159E9, 1.668666207E9, 1.668666255E9, 1.668666303E9, 1.668666351E9, 1.668666399E9, 1.668666447E9, 1.668666495E9, 1.668666543E9, 1.668666591E9, 1.668666639E9, 1.668666687E9, 1.668666735E9, 1.668666783E9, 1.668666831E9, 1.668666879E9, 1.668666927E9, 1.668666975E9, 1.668667023E9, 1.668667071E9, 1.668667119E9, 1.668667167E9, 1.668667215E9, 1.668667263E9, 1.668667311E9, 1.668667359E9, 1.668667407E9, 1.668667455E9, 1.668667503E9, 1.668667551E9, 1.668667599E9, 1.66866786E9, 1.66866804E9, 1.668673923E9, 1.668673971E9, 1.668674019E9, 1.668674067E9, 1.668674115E9, 1.668674163E9, 1.668674211E9, 1.668674259E9, 1.668674307E9, 1.668674355E9, 1.668674403E9, 1.668674451E9, 1.668674499E9, 1.668674547E9, 1.668674595E9, 1.668674643E9, 1.668674691E9, 1.668674739E9, 1.668674787E9, 1.668674835E9, 1.668674883E9, 1.668674931E9, 1.668674979E9, 1.668675027E9, 1.668675075E9, 1.668675123E9, 1.668675171E9, 1.668675219E9, 1.668675267E9, 1.668675315E9, 1.668675363E9, 1.668675411E9, 1.668675459E9, 1.668675507E9, 1.668675555E9, 1.668675603E9, 1.668675651E9, 1.668675699E9, 1.668675747E9, 1.668675795E9, 1.668675843E9, 1.668675891E9, 1.668675939E9, 1.668675987E9, 1.668676035E9, 1.668676083E9, 1.668676131E9, 1.668676179E9, 1.668676227E9, 1.668676275E9, 1.668676323E9, 1.668676371E9, 1.668676419E9, 1.668676467E9, 1.668676515E9, 1.668676563E9, 1.668676611E9, 1.668676659E9, 1.668676707E9, 1.668676755E9, 1.668676803E9, 1.668676851E9, 1.668676899E9, 1.668676947E9, 1.668676995E9, 1.668677043E9, 1.668677091E9, 1.668677139E9, 1.668677187E9, 1.668677235E9, 1.668677283E9, 1.668677331E9, 1.668677379E9, 1.6686777E9, 1.66867788E9, 1.668683621E9, 1.668683669E9, 1.668683717E9, 1.668683765E9, 1.668683813E9, 1.668683861E9, 1.668683909E9, 1.668683957E9, 1.668684005E9, 1.668684053E9, 1.668684101E9, 1.668684149E9, 1.668684197E9, 1.668684245E9, 1.668684293E9, 1.668684341E9, 1.668684389E9, 1.668684437E9, 1.668684485E9, 1.668684533E9, 1.668684581E9, 1.668684629E9, 1.668684677E9, 1.668684725E9, 1.668684773E9, 1.668684821E9, 1.668684869E9, 1.668684917E9, 1.668684965E9, 1.668685013E9, 1.668685061E9, 1.668685109E9, 1.668685157E9, 1.668685205E9, 1.668685253E9, 1.668685301E9, 1.668685349E9, 1.668685397E9, 1.668685445E9, 1.668685493E9, 1.668685541E9, 1.668685589E9, 1.668685637E9, 1.668685685E9, 1.668685733E9, 1.668685781E9, 1.668685829E9, 1.668685877E9, 1.668685925E9, 1.668685973E9, 1.668686021E9, 1.668686069E9, 1.668686117E9, 1.668686165E9, 1.668686213E9, 1.668686261E9, 1.668686309E9, 1.668686357E9, 1.668686405E9, 1.668686453E9, 1.668686501E9, 1.668686549E9, 1.668686597E9, 1.668686645E9, 1.668686693E9, 1.668686741E9, 1.668686789E9, 1.668686837E9, 1.668686885E9, 1.668686933E9, 1.668686981E9, 1.668687029E9, 1.66868742E9, 1.6686876E9, 1.668693376E9, 1.668693424E9, 1.668693472E9, 1.66869352E9, 1.668693568E9, 1.668693616E9, 1.668693664E9, 1.668693712E9, 1.66869376E9, 1.668693808E9, 1.668693856E9, 1.668693904E9, 1.668693952E9, 1.668694E9, 1.668694048E9, 1.668694096E9, 1.668694144E9, 1.668694192E9, 1.66869424E9, 1.668694288E9, 1.668694336E9, 1.668694384E9, 1.668694432E9, 1.66869448E9, 1.668694528E9, 1.668694576E9, 1.668694624E9, 1.668694672E9, 1.66869472E9, 1.668694768E9, 1.668694816E9, 1.668694864E9, 1.668694912E9, 1.66869496E9, 1.668695008E9, 1.668695056E9, 1.668695104E9, 1.668695152E9, 1.6686952E9, 1.668695248E9, 1.668695296E9, 1.668695344E9, 1.668695392E9, 1.66869544E9, 1.668695488E9, 1.668695536E9, 1.668695584E9, 1.668695632E9, 1.66869568E9, 1.668695728E9, 1.668695776E9, 1.668695824E9, 1.668695872E9, 1.66869592E9, 1.668695968E9, 1.668696016E9, 1.668696064E9, 1.668696112E9, 1.66869616E9, 1.668696208E9, 1.668696256E9, 1.668696304E9, 1.668696352E9, 1.6686964E9, 1.668696448E9, 1.668696496E9, 1.668696544E9, 1.668696592E9, 1.66869664E9, 1.668696688E9, 1.668696736E9, 1.668696784E9, 1.668696832E9, 1.66869688E9, 1.6686972E9, 1.66869738E9, 1.668703111E9, 1.668703159E9, 1.668703207E9, 1.668703255E9, 1.668703303E9, 1.668703351E9, 1.668703399E9, 1.668703447E9, 1.668703495E9, 1.668703543E9, 1.668703591E9, 1.668703639E9, 1.668703687E9, 1.668703735E9, 1.668703783E9, 1.668703831E9, 1.668703879E9, 1.668703927E9, 1.668703975E9, 1.668704023E9, 1.668704071E9, 1.668704119E9, 1.668704167E9, 1.668704215E9, 1.668704263E9, 1.668704311E9, 1.668704359E9, 1.668704407E9, 1.668704455E9, 1.668704503E9, 1.668704551E9, 1.668704599E9, 1.668704647E9, 1.668704695E9, 1.668704743E9, 1.668704791E9, 1.668704839E9, 1.668704887E9, 1.668704935E9, 1.668704983E9, 1.668705031E9, 1.668705079E9, 1.668705127E9, 1.668705175E9, 1.668705223E9, 1.668705271E9, 1.668705319E9, 1.668705367E9, 1.668705415E9, 1.668705463E9, 1.668705511E9, 1.668705559E9, 1.668705607E9, 1.668705655E9, 1.668705703E9, 1.668705751E9, 1.668705799E9, 1.668705847E9, 1.668705895E9, 1.668705943E9, 1.668705991E9, 1.668706039E9, 1.668706087E9, 1.668706135E9, 1.668706183E9, 1.668706231E9, 1.668706279E9, 1.668706327E9, 1.668706375E9, 1.668706423E9, 1.668706471E9, 1.668706519E9, 1.66870686E9, 1.66870704E9, 1.668712787E9, 1.668712835E9, 1.668712883E9, 1.668712931E9, 1.668712979E9, 1.668713027E9, 1.668713075E9, 1.668713123E9, 1.668713171E9, 1.668713219E9, 1.668713267E9, 1.668713315E9, 1.668713363E9, 1.668713411E9, 1.668713459E9, 1.668713507E9, 1.668713555E9, 1.668713603E9, 1.668713651E9, 1.668713699E9, 1.668713747E9, 1.668713795E9, 1.668713843E9, 1.668713891E9, 1.668713939E9, 1.668713987E9, 1.668714035E9, 1.668714083E9, 1.668714131E9, 1.668714179E9, 1.668714227E9, 1.668714275E9, 1.668714323E9, 1.668714371E9, 1.668714419E9, 1.668714467E9, 1.668714515E9, 1.668714563E9, 1.668714611E9, 1.668714659E9, 1.668714707E9, 1.668714755E9, 1.668714803E9, 1.668714851E9, 1.668714899E9, 1.668714947E9, 1.668714995E9, 1.668715043E9, 1.668715091E9, 1.668715139E9, 1.668715187E9, 1.668715235E9, 1.668715283E9, 1.668715331E9, 1.668715379E9, 1.668715427E9, 1.668715475E9, 1.668715523E9, 1.668715571E9, 1.668715619E9, 1.668715667E9, 1.668715715E9, 1.668715763E9, 1.668715811E9, 1.668715859E9, 1.668715907E9, 1.668715955E9, 1.668716003E9, 1.668716051E9, 1.668716099E9, 1.66871646E9, 1.66871664E9, 1.668722338E9, 1.668722386E9, 1.668722434E9, 1.668722482E9, 1.66872253E9, 1.668722578E9, 1.668722626E9, 1.668722674E9, 1.668722722E9, 1.66872277E9, 1.668722818E9, 1.668722866E9, 1.668722914E9, 1.668722962E9, 1.66872301E9, 1.668723058E9, 1.668723106E9, 1.668723154E9, 1.668723202E9, 1.66872325E9, 1.668723298E9, 1.668723346E9, 1.668723394E9, 1.668723442E9, 1.66872349E9, 1.668723538E9, 1.668723586E9, 1.668723634E9, 1.668723682E9, 1.66872373E9, 1.668723778E9, 1.668723826E9, 1.668723874E9, 1.668723922E9, 1.66872397E9, 1.668724018E9, 1.668724066E9, 1.668724114E9, 1.668724162E9, 1.66872421E9, 1.668724258E9, 1.668724306E9, 1.668724354E9, 1.668724402E9, 1.66872445E9, 1.668724498E9, 1.668724546E9, 1.668724594E9, 1.668724642E9, 1.66872469E9, 1.668724738E9, 1.668724786E9, 1.668724834E9, 1.668724882E9, 1.66872493E9, 1.668724978E9, 1.668725026E9, 1.668725074E9, 1.668725122E9, 1.66872517E9, 1.668725218E9, 1.668725266E9, 1.668725314E9, 1.668725362E9, 1.66872541E9, 1.668725458E9, 1.668725506E9, 1.668725554E9, 1.668725602E9, 1.66872565E9, 1.668726E9, 1.66872618E9, 1.668731894E9, 1.668731942E9, 1.66873199E9, 1.668732038E9, 1.668732086E9, 1.668732134E9, 1.668732182E9, 1.66873223E9, 1.668732278E9, 1.668732326E9, 1.668732374E9, 1.668732422E9, 1.66873247E9, 1.668732518E9, 1.668732566E9, 1.668732614E9, 1.668732662E9, 1.66873271E9, 1.668732758E9, 1.668732806E9, 1.668732854E9, 1.668732902E9, 1.66873295E9, 1.668732998E9, 1.668733046E9, 1.668733094E9, 1.668733142E9, 1.66873319E9, 1.668733238E9, 1.668733286E9, 1.668733334E9, 1.668733382E9, 1.66873343E9, 1.668733478E9, 1.668733526E9, 1.668733574E9, 1.668733622E9, 1.66873367E9, 1.668733718E9, 1.668733766E9, 1.668733814E9, 1.668733862E9, 1.66873391E9, 1.668733958E9, 1.668734006E9, 1.668734054E9, 1.668734102E9, 1.66873415E9, 1.668734198E9, 1.668734246E9, 1.668734294E9, 1.668734342E9, 1.66873439E9, 1.668734438E9, 1.668734486E9, 1.668734534E9, 1.668734582E9, 1.66873463E9, 1.668734678E9, 1.668734726E9, 1.668734774E9, 1.668734822E9, 1.66873487E9, 1.668734918E9, 1.668734966E9, 1.668735014E9, 1.668735062E9, 1.66873511E9, 1.668735158E9, 1.668735206E9, 1.668735254E9, 1.668735302E9, 1.66873535E9, 1.6687356E9, 1.66873578E9, 1.66874151E9, 1.668741558E9, 1.668741606E9, 1.668741654E9, 1.668741702E9, 1.66874175E9, 1.668741798E9, 1.668741846E9, 1.668741894E9, 1.668741942E9, 1.66874199E9, 1.668742038E9, 1.668742086E9, 1.668742134E9, 1.668742182E9, 1.66874223E9, 1.668742278E9, 1.668742326E9, 1.668742374E9, 1.668742422E9, 1.66874247E9, 1.668742518E9, 1.668742566E9, 1.668742614E9, 1.668742662E9, 1.66874271E9, 1.668742758E9, 1.668742806E9, 1.668742854E9, 1.668742902E9, 1.66874295E9, 1.668742998E9, 1.668743046E9, 1.668743094E9, 1.668743142E9, 1.66874319E9, 1.668743238E9, 1.668743286E9, 1.668743334E9, 1.668743382E9, 1.66874343E9, 1.668743478E9, 1.668743526E9, 1.668743574E9, 1.668743622E9, 1.66874367E9, 1.668743718E9, 1.668743766E9, 1.668743814E9, 1.668743862E9, 1.66874391E9, 1.668743958E9, 1.668744006E9, 1.668744054E9, 1.668744102E9, 1.66874415E9, 1.668744198E9, 1.668744246E9, 1.668744294E9, 1.668744342E9, 1.66874439E9, 1.668744438E9, 1.668744486E9, 1.668744534E9, 1.668744582E9, 1.66874463E9, 1.668744678E9, 1.668744726E9, 1.668744774E9, 1.668744822E9, 1.66874487E9, 1.66874526E9, 1.66874544E9, 1.66875103E9, 1.668751078E9, 1.668751126E9, 1.668751174E9, 1.668751222E9, 1.66875127E9, 1.668751318E9, 1.668751366E9, 1.668751414E9, 1.668751462E9, 1.66875151E9, 1.668751558E9, 1.668751606E9, 1.668751654E9, 1.668751702E9, 1.66875175E9, 1.668751798E9, 1.668751846E9, 1.668751894E9, 1.668751942E9, 1.66875199E9, 1.668752038E9, 1.668752086E9, 1.668752134E9, 1.668752182E9, 1.66875223E9, 1.668752278E9, 1.668752326E9, 1.668752374E9, 1.668752422E9, 1.66875247E9, 1.668752518E9, 1.668752566E9, 1.668752614E9, 1.668752662E9, 1.66875271E9, 1.668752758E9, 1.668752806E9, 1.668752854E9, 1.668752902E9, 1.66875295E9, 1.668752998E9, 1.668753046E9, 1.668753094E9, 1.668753142E9, 1.66875319E9, 1.668753238E9, 1.668753286E9, 1.668753334E9, 1.668753382E9, 1.66875343E9, 1.668753478E9, 1.668753526E9, 1.668753574E9, 1.668753622E9, 1.66875367E9, 1.668753718E9, 1.668753766E9, 1.668753814E9, 1.668753862E9, 1.66875391E9, 1.668753958E9, 1.668754006E9, 1.668754054E9, 1.668754102E9, 1.66875415E9, 1.668754198E9, 1.668754246E9, 1.668754294E9, 1.668754342E9, 1.66875439E9, 1.66875468E9, 1.66875486E9, 1.668760559E9, 1.668760607E9, 1.668760655E9, 1.668760703E9, 1.668760751E9, 1.668760799E9, 1.668760847E9, 1.668760895E9, 1.668760943E9, 1.668760991E9, 1.668761039E9, 1.668761087E9, 1.668761135E9, 1.668761183E9, 1.668761231E9, 1.668761279E9, 1.668761327E9, 1.668761375E9, 1.668761423E9, 1.668761471E9, 1.668761519E9, 1.668761567E9, 1.668761615E9, 1.668761663E9, 1.668761711E9, 1.668761759E9, 1.668761807E9, 1.668761855E9, 1.668761903E9, 1.668761951E9, 1.668761999E9, 1.668762047E9, 1.668762095E9, 1.668762143E9, 1.668762191E9, 1.668762239E9, 1.668762287E9, 1.668762335E9, 1.668762383E9, 1.668762431E9, 1.668762479E9, 1.668762527E9, 1.668762575E9, 1.668762623E9, 1.668762671E9, 1.668762719E9, 1.668762767E9, 1.668762815E9, 1.668762863E9, 1.668762911E9, 1.668762959E9, 1.668763007E9, 1.668763055E9, 1.668763103E9, 1.668763151E9, 1.668763199E9, 1.668763247E9, 1.668763295E9, 1.668763343E9, 1.668763391E9, 1.668763439E9, 1.668763487E9, 1.668763535E9, 1.668763583E9, 1.668763631E9, 1.668763679E9, 1.668763727E9, 1.668763775E9, 1.668763823E9, 1.668763871E9, 1.668763919E9, 1.66876422E9, 1.6687644E9, 1.668770084E9, 1.668770132E9, 1.66877018E9, 1.668770228E9, 1.668770276E9, 1.668770324E9, 1.668770372E9, 1.66877042E9, 1.668770468E9, 1.668770516E9, 1.668770564E9, 1.668770612E9, 1.66877066E9, 1.668770708E9, 1.668770756E9, 1.668770804E9, 1.668770852E9, 1.6687709E9, 1.668770948E9, 1.668770996E9, 1.668771044E9, 1.668771092E9, 1.66877114E9, 1.668771188E9, 1.668771236E9, 1.668771284E9, 1.668771332E9, 1.66877138E9, 1.668771428E9, 1.668771476E9, 1.668771524E9, 1.668771572E9, 1.66877162E9, 1.668771668E9, 1.668771716E9, 1.668771764E9, 1.668771812E9, 1.66877186E9, 1.668771908E9, 1.668771956E9, 1.668772004E9, 1.668772052E9, 1.6687721E9, 1.668772148E9, 1.668772196E9, 1.668772244E9, 1.668772292E9, 1.66877234E9, 1.668772388E9, 1.668772436E9, 1.668772484E9, 1.668772532E9, 1.66877258E9, 1.668772628E9, 1.668772676E9, 1.668772724E9, 1.668772772E9, 1.66877282E9, 1.668772868E9, 1.668772916E9, 1.668772964E9, 1.668773012E9, 1.66877306E9, 1.668773108E9, 1.668773156E9, 1.668773204E9, 1.668773252E9, 1.6687733E9, 1.668773348E9, 1.668773396E9, 1.668773444E9, 1.668773492E9, 1.66877354E9, 1.66877394E9, 1.66877412E9, 1.668780077E9, 1.668780125E9, 1.668780173E9, 1.668780221E9, 1.668780269E9, 1.668780317E9, 1.668780365E9, 1.668780413E9, 1.668780461E9, 1.668780509E9, 1.668780557E9, 1.668780605E9, 1.668780653E9, 1.668780701E9, 1.668780749E9, 1.668780797E9, 1.668780845E9, 1.668780893E9, 1.668780941E9, 1.668780989E9, 1.668781037E9, 1.668781085E9, 1.668781133E9, 1.668781181E9, 1.668781229E9, 1.668781277E9, 1.668781325E9, 1.668781373E9, 1.668781421E9, 1.668781469E9, 1.668781517E9, 1.668781565E9, 1.668781613E9, 1.668781661E9, 1.668781709E9, 1.668781757E9, 1.668781805E9, 1.668781853E9, 1.668781901E9, 1.668781949E9, 1.668781997E9, 1.668782045E9, 1.668782093E9, 1.668782141E9, 1.668782189E9, 1.668782237E9, 1.668782285E9, 1.668782333E9, 1.668782381E9, 1.668782429E9, 1.668782477E9, 1.668782525E9, 1.668782573E9, 1.668782621E9, 1.668782669E9, 1.668782717E9, 1.668782765E9, 1.668782813E9, 1.668782861E9, 1.668782909E9, 1.668782957E9, 1.668783005E9, 1.668783053E9, 1.668783101E9, 1.668783149E9, 1.668783197E9, 1.668783245E9, 1.668783293E9, 1.668783341E9, 1.668783389E9, 1.66878378E9, 1.668783781E9, 1.668789398E9, 1.668789446E9, 1.668789494E9, 1.668789542E9, 1.66878959E9, 1.668789638E9, 1.668789686E9, 1.668789734E9, 1.668789782E9, 1.66878983E9, 1.668789878E9, 1.668789926E9, 1.668789974E9, 1.668790022E9, 1.66879007E9, 1.668790118E9, 1.668790166E9, 1.668790214E9, 1.668790262E9, 1.66879031E9, 1.668790358E9, 1.668790406E9, 1.668790454E9, 1.668790502E9, 1.66879055E9, 1.668790598E9, 1.668790646E9, 1.668790694E9, 1.668790742E9, 1.66879079E9, 1.668790838E9, 1.668790886E9, 1.668790934E9, 1.668790982E9, 1.66879103E9, 1.668791078E9, 1.668791126E9, 1.668791174E9, 1.668791222E9, 1.66879127E9, 1.668791318E9, 1.668791366E9, 1.668791414E9, 1.668791462E9, 1.66879151E9, 1.668791558E9, 1.668791606E9, 1.668791654E9, 1.668791702E9, 1.66879175E9, 1.668791798E9, 1.668791846E9, 1.668791894E9, 1.668791942E9, 1.66879199E9, 1.668792038E9, 1.668792086E9, 1.668792134E9, 1.668792182E9, 1.66879223E9, 1.668792278E9, 1.668792326E9, 1.668792374E9, 1.668792422E9, 1.66879247E9, 1.668792518E9, 1.668792566E9, 1.668792614E9, 1.668792662E9, 1.66879271E9, 1.66879302E9, 1.6687932E9, 1.668798926E9, 1.668798974E9, 1.668799022E9, 1.66879907E9, 1.668799118E9, 1.668799166E9, 1.668799214E9, 1.668799262E9, 1.66879931E9, 1.668799358E9, 1.668799406E9, 1.668799454E9, 1.668799502E9, 1.66879955E9, 1.668799598E9, 1.668799646E9, 1.668799694E9, 1.668799742E9, 1.66879979E9, 1.668799838E9, 1.668799886E9, 1.668799934E9, 1.668799982E9, 1.66880003E9, 1.668800078E9, 1.668800126E9, 1.668800174E9, 1.668800222E9, 1.66880027E9, 1.668800318E9, 1.668800366E9, 1.668800414E9, 1.668800462E9, 1.66880051E9, 1.668800558E9, 1.668800606E9, 1.668800654E9, 1.668800702E9, 1.66880075E9, 1.668800798E9, 1.668800846E9, 1.668800894E9, 1.668800942E9, 1.66880099E9, 1.668801038E9, 1.668801086E9, 1.668801134E9, 1.668801182E9, 1.66880123E9, 1.668801278E9, 1.668801326E9, 1.668801374E9, 1.668801422E9, 1.66880147E9, 1.668801518E9, 1.668801566E9, 1.668801614E9, 1.668801662E9, 1.66880171E9, 1.668801758E9, 1.668801806E9, 1.668801854E9, 1.668801902E9, 1.66880195E9, 1.668801998E9, 1.668802046E9, 1.668802094E9, 1.668802142E9, 1.66880219E9, 1.668802238E9, 1.668802286E9, 1.668802334E9, 1.668802382E9, 1.66880243E9, 1.6688028E9, 1.66880298E9, 1.668808649E9, 1.668808697E9, 1.668808745E9, 1.668808793E9, 1.668808841E9, 1.668808889E9, 1.668808937E9, 1.668808985E9, 1.668809033E9, 1.668809081E9, 1.668809129E9, 1.668809177E9, 1.668809225E9, 1.668809273E9, 1.668809321E9, 1.668809369E9, 1.668809417E9, 1.668809465E9, 1.668809513E9, 1.668809561E9, 1.668809609E9, 1.668809657E9, 1.668809705E9, 1.668809753E9, 1.668809801E9, 1.668809849E9, 1.668809897E9, 1.668809945E9, 1.668809993E9, 1.668810041E9, 1.668810089E9, 1.668810137E9, 1.668810185E9, 1.668810233E9, 1.668810281E9, 1.668810329E9, 1.668810377E9, 1.668810425E9, 1.668810473E9, 1.668810521E9, 1.668810569E9, 1.668810617E9, 1.668810665E9, 1.668810713E9, 1.668810761E9, 1.668810809E9, 1.668810857E9, 1.668810905E9, 1.668810953E9, 1.668811001E9, 1.668811049E9, 1.668811097E9, 1.668811145E9, 1.668811193E9, 1.668811241E9, 1.668811289E9, 1.668811337E9, 1.668811385E9, 1.668811433E9, 1.668811481E9, 1.668811529E9, 1.668811577E9, 1.668811625E9, 1.668811673E9, 1.668811721E9, 1.668811769E9, 1.668811817E9, 1.668811865E9, 1.668811913E9, 1.668811961E9, 1.668812009E9, 1.66881234E9, 1.66881252E9, 1.668818342E9, 1.66881839E9, 1.668818438E9, 1.668818486E9, 1.668818534E9, 1.668818582E9, 1.66881863E9, 1.668818678E9, 1.668818726E9, 1.668818774E9, 1.668818822E9, 1.66881887E9, 1.668818918E9, 1.668818966E9, 1.668819014E9, 1.668819062E9, 1.66881911E9, 1.668819158E9, 1.668819206E9, 1.668819254E9, 1.668819302E9, 1.66881935E9, 1.668819398E9, 1.668819446E9, 1.668819494E9, 1.668819542E9, 1.66881959E9, 1.668819638E9, 1.668819686E9, 1.668819734E9, 1.668819782E9, 1.66881983E9, 1.668819878E9, 1.668819926E9, 1.668819974E9, 1.668820022E9, 1.66882007E9, 1.668820118E9, 1.668820166E9, 1.668820214E9, 1.668820262E9, 1.66882031E9, 1.668820358E9, 1.668820406E9, 1.668820454E9, 1.668820502E9, 1.66882055E9, 1.668820598E9, 1.668820646E9, 1.668820694E9, 1.668820742E9, 1.66882079E9, 1.668820838E9, 1.668820886E9, 1.668820934E9, 1.668820982E9, 1.66882103E9, 1.668821078E9, 1.668821126E9, 1.668821174E9, 1.668821222E9, 1.66882127E9, 1.668821318E9, 1.668821366E9, 1.668821414E9, 1.668821462E9, 1.66882151E9, 1.668821558E9, 1.668821606E9, 1.668821654E9, 1.668821702E9, 1.66882175E9, 1.668822E9, 1.66882218E9, 1.668827872E9, 1.66882792E9, 1.668827968E9, 1.668828016E9, 1.668828064E9, 1.668828112E9, 1.66882816E9, 1.668828208E9, 1.668828256E9, 1.668828304E9, 1.668828352E9, 1.6688284E9, 1.668828448E9, 1.668828496E9, 1.668828544E9, 1.668828592E9, 1.66882864E9, 1.668828688E9, 1.668828736E9, 1.668828784E9, 1.668828832E9, 1.66882888E9, 1.668828928E9, 1.668828976E9, 1.668829024E9, 1.668829072E9, 1.66882912E9, 1.668829168E9, 1.668829216E9, 1.668829264E9, 1.668829312E9, 1.66882936E9, 1.668829408E9, 1.668829456E9, 1.668829504E9, 1.668829552E9, 1.6688296E9, 1.668829648E9, 1.668829696E9, 1.668829744E9, 1.668829792E9, 1.66882984E9, 1.668829888E9, 1.668829936E9, 1.668829984E9, 1.668830032E9, 1.66883008E9, 1.668830128E9, 1.668830176E9, 1.668830224E9, 1.668830272E9, 1.66883032E9, 1.668830368E9, 1.668830416E9, 1.668830464E9, 1.668830512E9, 1.66883056E9, 1.668830608E9, 1.668830656E9, 1.668830704E9, 1.668830752E9, 1.6688308E9, 1.668830848E9, 1.668830896E9, 1.668830944E9, 1.668830992E9, 1.66883104E9, 1.668831088E9, 1.668831136E9, 1.668831184E9, 1.668831232E9, 1.66883128E9, 1.66883166E9, 1.66883184E9, 1.66883755E9, 1.668837598E9, 1.668837646E9, 1.668837694E9, 1.668837742E9, 1.66883779E9, 1.668837838E9, 1.668837886E9, 1.668837934E9, 1.668837982E9, 1.66883803E9, 1.668838078E9, 1.668838126E9, 1.668838174E9, 1.668838222E9, 1.66883827E9, 1.668838318E9, 1.668838366E9, 1.668838414E9, 1.668838462E9, 1.66883851E9, 1.668838558E9, 1.668838606E9, 1.668838654E9, 1.668838702E9, 1.66883875E9, 1.668838798E9, 1.668838846E9, 1.668838894E9, 1.668838942E9, 1.66883899E9, 1.668839038E9, 1.668839086E9, 1.668839134E9, 1.668839182E9, 1.66883923E9, 1.668839278E9, 1.668839326E9, 1.668839374E9, 1.668839422E9, 1.66883947E9, 1.668839518E9, 1.668839566E9, 1.668839614E9, 1.668839662E9, 1.66883971E9, 1.668839758E9, 1.668839806E9, 1.668839854E9, 1.668839902E9, 1.66883995E9, 1.668839998E9, 1.668840046E9, 1.668840094E9, 1.668840142E9, 1.66884019E9, 1.668840238E9, 1.668840286E9, 1.668840334E9, 1.668840382E9, 1.66884043E9, 1.668840478E9, 1.668840526E9, 1.668840574E9, 1.668840622E9, 1.66884067E9, 1.668840718E9, 1.668840766E9, 1.668840814E9, 1.668840862E9, 1.66884091E9, 1.66884126E9, 1.66884144E9, 1.668847184E9, 1.668847232E9, 1.66884728E9, 1.668847328E9, 1.668847376E9, 1.668847424E9, 1.668847472E9, 1.66884752E9, 1.668847568E9, 1.668847616E9, 1.668847664E9, 1.668847712E9, 1.66884776E9, 1.668847808E9, 1.668847856E9, 1.668847904E9, 1.668847952E9, 1.668848E9, 1.668848048E9, 1.668848096E9, 1.668848144E9, 1.668848192E9, 1.66884824E9, 1.668848288E9, 1.668848336E9, 1.668848384E9, 1.668848432E9, 1.66884848E9, 1.668848528E9, 1.668848576E9, 1.668848624E9, 1.668848672E9, 1.66884872E9, 1.668848768E9, 1.668848816E9, 1.668848864E9, 1.668848912E9, 1.66884896E9, 1.668849008E9, 1.668849056E9, 1.668849104E9, 1.668849152E9, 1.6688492E9, 1.668849248E9, 1.668849296E9, 1.668849344E9, 1.668849392E9, 1.66884944E9, 1.668849488E9, 1.668849536E9, 1.668849584E9, 1.668849632E9, 1.66884968E9, 1.668849728E9, 1.668849776E9, 1.668849824E9, 1.668849872E9, 1.66884992E9, 1.668849968E9, 1.668850016E9, 1.668850064E9, 1.668850112E9, 1.66885016E9, 1.668850208E9, 1.668850256E9, 1.668850304E9, 1.668850352E9, 1.6688504E9, 1.668850448E9, 1.668850496E9, 1.668850544E9, 1.668850592E9, 1.66885064E9, 1.66885092E9, 1.66885116E9, 1.668856948E9, 1.668856996E9, 1.668857044E9, 1.668857092E9, 1.66885714E9, 1.668857188E9, 1.668857236E9, 1.668857284E9, 1.668857332E9, 1.66885738E9, 1.668857428E9, 1.668857476E9, 1.668857524E9, 1.668857572E9, 1.66885762E9, 1.668857668E9, 1.668857716E9, 1.668857764E9, 1.668857812E9, 1.66885786E9, 1.668857908E9, 1.668857956E9, 1.668858004E9, 1.668858052E9, 1.6688581E9, 1.668858148E9, 1.668858196E9, 1.668858244E9, 1.668858292E9, 1.66885834E9, 1.668858388E9, 1.668858436E9, 1.668858484E9, 1.668858532E9, 1.66885858E9, 1.668858628E9, 1.668858676E9, 1.668858724E9, 1.668858772E9, 1.66885882E9, 1.668858868E9, 1.668858916E9, 1.668858964E9, 1.668859012E9, 1.66885906E9, 1.668859108E9, 1.668859156E9, 1.668859204E9, 1.668859252E9, 1.6688593E9, 1.668859348E9, 1.668859396E9, 1.668859444E9, 1.668859492E9, 1.66885954E9, 1.668859588E9, 1.668859636E9, 1.668859684E9, 1.668859732E9, 1.66885978E9, 1.668859828E9, 1.668859876E9, 1.668859924E9, 1.668859972E9, 1.66886002E9, 1.668860068E9, 1.668860116E9, 1.668860164E9, 1.668860212E9, 1.66886026E9, 1.66886064E9, 1.66886082E9, 1.668866924E9, 1.668866972E9, 1.66886702E9, 1.668867068E9, 1.668867116E9, 1.668867164E9, 1.668867212E9, 1.66886726E9, 1.668867308E9, 1.668867356E9, 1.668867404E9, 1.668867452E9, 1.6688675E9, 1.668867548E9, 1.668867596E9, 1.668867644E9, 1.668867692E9, 1.66886774E9, 1.668867788E9, 1.668867836E9, 1.668867884E9, 1.668867932E9, 1.66886798E9, 1.668868028E9, 1.668868076E9, 1.668868124E9, 1.668868172E9, 1.66886822E9, 1.668868268E9, 1.668868316E9, 1.668868364E9, 1.668868412E9, 1.66886846E9, 1.668868508E9, 1.668868556E9, 1.668868604E9, 1.668868652E9, 1.6688687E9, 1.668868748E9, 1.668868796E9, 1.668868844E9, 1.668868892E9, 1.66886894E9, 1.668868988E9, 1.668869036E9, 1.668869084E9, 1.668869132E9, 1.66886918E9, 1.668869228E9, 1.668869276E9, 1.668869324E9, 1.668869372E9, 1.66886942E9, 1.668869468E9, 1.668869516E9, 1.668869564E9, 1.668869612E9, 1.66886966E9, 1.668869708E9, 1.668869756E9, 1.668869804E9, 1.668869852E9, 1.6688699E9, 1.668869948E9, 1.668869996E9, 1.668870044E9, 1.668870092E9, 1.66887014E9, 1.668870188E9, 1.668870236E9, 1.668870284E9, 1.668870332E9, 1.66887038E9, 1.66887066E9, 1.66887084E9, 1.668876543E9, 1.668876591E9, 1.668876639E9, 1.668876687E9, 1.668876735E9, 1.668876783E9, 1.668876831E9, 1.668876879E9, 1.668876927E9, 1.668876975E9, 1.668877023E9, 1.668877071E9, 1.668877119E9, 1.668877167E9, 1.668877215E9, 1.668877263E9, 1.668877311E9, 1.668877359E9, 1.668877407E9, 1.668877455E9, 1.668877503E9, 1.668877551E9, 1.668877599E9, 1.668877647E9, 1.668877695E9, 1.668877743E9, 1.668877791E9, 1.668877839E9, 1.668877887E9, 1.668877935E9, 1.668877983E9, 1.668878031E9, 1.668878079E9, 1.668878127E9, 1.668878175E9, 1.668878223E9, 1.668878271E9, 1.668878319E9, 1.668878367E9, 1.668878415E9, 1.668878463E9, 1.668878511E9, 1.668878559E9, 1.668878607E9, 1.668878655E9, 1.668878703E9, 1.668878751E9, 1.668878799E9, 1.668878847E9, 1.668878895E9, 1.668878943E9, 1.668878991E9, 1.668879039E9, 1.668879087E9, 1.668879135E9, 1.668879183E9, 1.668879231E9, 1.668879279E9, 1.668879327E9, 1.668879375E9, 1.668879423E9, 1.668879471E9, 1.668879519E9, 1.668879567E9, 1.668879615E9, 1.668879663E9, 1.668879711E9, 1.668879759E9, 1.668879807E9, 1.668879855E9, 1.668879903E9, 1.668879951E9, 1.668879999E9, 1.66888032E9, 1.6688805E9, 1.668886185E9, 1.668886233E9, 1.668886281E9, 1.668886329E9, 1.668886377E9, 1.668886425E9, 1.668886473E9, 1.668886521E9, 1.668886569E9, 1.668886617E9, 1.668886665E9, 1.668886713E9, 1.668886761E9, 1.668886809E9, 1.668886857E9, 1.668886905E9, 1.668886953E9, 1.668887001E9, 1.668887049E9, 1.668887097E9, 1.668887145E9, 1.668887193E9, 1.668887241E9, 1.668887289E9, 1.668887337E9, 1.668887385E9, 1.668887433E9, 1.668887481E9, 1.668887529E9, 1.668887577E9, 1.668887625E9, 1.668887673E9, 1.668887721E9, 1.668887769E9, 1.668887817E9, 1.668887865E9, 1.668887913E9, 1.668887961E9, 1.668888009E9, 1.668888057E9, 1.668888105E9, 1.668888153E9, 1.668888201E9, 1.668888249E9, 1.668888297E9, 1.668888345E9, 1.668888393E9, 1.668888441E9, 1.668888489E9, 1.668888537E9, 1.668888585E9, 1.668888633E9, 1.668888681E9, 1.668888729E9, 1.668888777E9, 1.668888825E9, 1.668888873E9, 1.668888921E9, 1.668888969E9, 1.668889017E9, 1.668889065E9, 1.668889113E9, 1.668889161E9, 1.668889209E9, 1.668889257E9, 1.668889305E9, 1.668889353E9, 1.668889401E9, 1.668889449E9, 1.668889497E9, 1.668889545E9, 1.668889593E9, 1.668889641E9, 1.668889689E9, 1.66888998E9, 1.66889016E9, 1.668895859E9, 1.668895907E9, 1.668895955E9, 1.668896003E9, 1.668896051E9, 1.668896099E9, 1.668896147E9, 1.668896195E9, 1.668896243E9, 1.668896291E9, 1.668896339E9, 1.668896387E9, 1.668896435E9, 1.668896483E9, 1.668896531E9, 1.668896579E9, 1.668896627E9, 1.668896675E9, 1.668896723E9, 1.668896771E9, 1.668896819E9, 1.668896867E9, 1.668896915E9, 1.668896963E9, 1.668897011E9, 1.668897059E9, 1.668897107E9, 1.668897155E9, 1.668897203E9, 1.668897251E9, 1.668897299E9, 1.668897347E9, 1.668897395E9, 1.668897443E9, 1.668897491E9, 1.668897539E9, 1.668897587E9, 1.668897635E9, 1.668897683E9, 1.668897731E9, 1.668897779E9, 1.668897827E9, 1.668897875E9, 1.668897923E9, 1.668897971E9, 1.668898019E9, 1.668898067E9, 1.668898115E9, 1.668898163E9, 1.668898211E9, 1.668898259E9, 1.668898307E9, 1.668898355E9, 1.668898403E9, 1.668898451E9, 1.668898499E9, 1.668898547E9, 1.668898595E9, 1.668898643E9, 1.668898691E9, 1.668898739E9, 1.668898787E9, 1.668898835E9, 1.668898883E9, 1.668898931E9, 1.668898979E9, 1.668899027E9, 1.668899075E9, 1.668899123E9, 1.668899171E9, 1.668899219E9, 1.66889958E9, 1.6688997E9, 1.668905375E9, 1.668905423E9, 1.668905471E9, 1.668905519E9, 1.668905567E9, 1.668905615E9, 1.668905663E9, 1.668905711E9, 1.668905759E9, 1.668905807E9, 1.668905855E9, 1.668905903E9, 1.668905951E9, 1.668905999E9, 1.668906047E9, 1.668906095E9, 1.668906143E9, 1.668906191E9, 1.668906239E9, 1.668906287E9, 1.668906335E9, 1.668906383E9, 1.668906431E9, 1.668906479E9, 1.668906527E9, 1.668906575E9, 1.668906623E9, 1.668906671E9, 1.668906719E9, 1.668906767E9, 1.668906815E9, 1.668906863E9, 1.668906911E9, 1.668906959E9, 1.668907007E9, 1.668907055E9, 1.668907103E9, 1.668907151E9, 1.668907199E9, 1.668907247E9, 1.668907295E9, 1.668907343E9, 1.668907391E9, 1.668907439E9, 1.668907487E9, 1.668907535E9, 1.668907583E9, 1.668907631E9, 1.668907679E9, 1.668907727E9, 1.668907775E9, 1.668907823E9, 1.668907871E9, 1.668907919E9, 1.668907967E9, 1.668908015E9, 1.668908063E9, 1.668908111E9, 1.668908159E9, 1.668908207E9, 1.668908255E9, 1.668908303E9, 1.668908351E9, 1.668908399E9, 1.668908447E9, 1.668908495E9, 1.668908543E9, 1.668908591E9, 1.668908639E9, 1.668908687E9, 1.668908735E9, 1.668908783E9, 1.668908831E9, 1.668908879E9, 1.668908927E9, 1.668908975E9, 1.668909023E9, 1.668909071E9, 1.668909119E9, 1.66890936E9, 1.66890954E9, 1.668915359E9, 1.668915407E9, 1.668915455E9, 1.668915503E9, 1.668915551E9, 1.668915599E9, 1.668915647E9, 1.668915695E9, 1.668915743E9, 1.668915791E9, 1.668915839E9, 1.668915887E9, 1.668915935E9, 1.668915983E9, 1.668916031E9, 1.668916079E9, 1.668916127E9, 1.668916175E9, 1.668916223E9, 1.668916271E9, 1.668916319E9, 1.668916367E9, 1.668916415E9, 1.668916463E9, 1.668916511E9, 1.668916559E9, 1.668916607E9, 1.668916655E9, 1.668916703E9, 1.668916751E9, 1.668916799E9, 1.668916847E9, 1.668916895E9, 1.668916943E9, 1.668916991E9, 1.668917039E9, 1.668917087E9, 1.668917135E9, 1.668917183E9, 1.668917231E9, 1.668917279E9, 1.668917327E9, 1.668917375E9, 1.668917423E9, 1.668917471E9, 1.668917519E9, 1.668917567E9, 1.668917615E9, 1.668917663E9, 1.668917711E9, 1.668917759E9, 1.668917807E9, 1.668917855E9, 1.668917903E9, 1.668917951E9, 1.668917999E9, 1.668918047E9, 1.668918095E9, 1.668918143E9, 1.668918191E9, 1.668918239E9, 1.668918287E9, 1.668918335E9, 1.668918383E9, 1.668918431E9, 1.668918479E9, 1.668918527E9, 1.668918575E9, 1.668918623E9, 1.668918671E9, 1.668918719E9, 1.66891902E9, 1.6689192E9, 1.668924855E9, 1.668924903E9, 1.668924951E9, 1.668924999E9, 1.668925047E9, 1.668925095E9, 1.668925143E9, 1.668925191E9, 1.668925239E9, 1.668925287E9, 1.668925335E9, 1.668925383E9, 1.668925431E9, 1.668925479E9, 1.668925527E9, 1.668925575E9, 1.668925623E9, 1.668925671E9, 1.668925719E9, 1.668925767E9, 1.668925815E9, 1.668925863E9, 1.668925911E9, 1.668925959E9, 1.668926007E9, 1.668926055E9, 1.668926103E9, 1.668926151E9, 1.668926199E9, 1.668926247E9, 1.668926295E9, 1.668926343E9, 1.668926391E9, 1.668926439E9, 1.668926487E9, 1.668926535E9, 1.668926583E9, 1.668926631E9, 1.668926679E9, 1.668926727E9, 1.668926775E9, 1.668926823E9, 1.668926871E9, 1.668926919E9, 1.668926967E9, 1.668927015E9, 1.668927063E9, 1.668927111E9, 1.668927159E9, 1.668927207E9, 1.668927255E9, 1.668927303E9, 1.668927351E9, 1.668927399E9, 1.668927447E9, 1.668927495E9, 1.668927543E9, 1.668927591E9, 1.668927639E9, 1.668927687E9, 1.668927735E9, 1.668927783E9, 1.668927831E9, 1.668927879E9, 1.668927927E9, 1.668927975E9, 1.668928023E9, 1.668928071E9, 1.668928119E9, 1.668928167E9, 1.668928215E9, 1.668928263E9, 1.668928311E9, 1.668928359E9, 1.66892862E9, 1.6689288E9, 1.668934503E9, 1.668934551E9, 1.668934599E9, 1.668934647E9, 1.668934695E9, 1.668934743E9, 1.668934791E9, 1.668934839E9, 1.668934887E9, 1.668934935E9, 1.668934983E9, 1.668935031E9, 1.668935079E9, 1.668935127E9, 1.668935175E9, 1.668935223E9, 1.668935271E9, 1.668935319E9, 1.668935367E9, 1.668935415E9, 1.668935463E9, 1.668935511E9, 1.668935559E9, 1.668935607E9, 1.668935655E9, 1.668935703E9, 1.668935751E9, 1.668935799E9, 1.668935847E9, 1.668935895E9, 1.668935943E9, 1.668935991E9, 1.668936039E9, 1.668936087E9, 1.668936135E9, 1.668936183E9, 1.668936231E9, 1.668936279E9, 1.668936327E9, 1.668936375E9, 1.668936423E9, 1.668936471E9, 1.668936519E9, 1.668936567E9, 1.668936615E9, 1.668936663E9, 1.668936711E9, 1.668936759E9, 1.668936807E9, 1.668936855E9, 1.668936903E9, 1.668936951E9, 1.668936999E9, 1.668937047E9, 1.668937095E9, 1.668937143E9, 1.668937191E9, 1.668937239E9, 1.668937287E9, 1.668937335E9, 1.668937383E9, 1.668937431E9, 1.668937479E9, 1.668937527E9, 1.668937575E9, 1.668937623E9, 1.668937671E9, 1.668937719E9, 1.668937767E9, 1.668937815E9, 1.668937863E9, 1.668937911E9, 1.668937959E9, 1.66893822E9, 1.66893846E9, 1.668944184E9, 1.668944232E9, 1.66894428E9, 1.668944328E9, 1.668944376E9, 1.668944424E9, 1.668944472E9, 1.66894452E9, 1.668944568E9, 1.668944616E9, 1.668944664E9, 1.668944712E9, 1.66894476E9, 1.668944808E9, 1.668944856E9, 1.668944904E9, 1.668944952E9, 1.668945E9, 1.668945048E9, 1.668945096E9, 1.668945144E9, 1.668945192E9, 1.66894524E9, 1.668945288E9, 1.668945336E9, 1.668945384E9, 1.668945432E9, 1.66894548E9, 1.668945528E9, 1.668945576E9, 1.668945624E9, 1.668945672E9, 1.66894572E9, 1.668945768E9, 1.668945816E9, 1.668945864E9, 1.668945912E9, 1.66894596E9, 1.668946008E9, 1.668946056E9, 1.668946104E9, 1.668946152E9, 1.6689462E9, 1.668946248E9, 1.668946296E9, 1.668946344E9, 1.668946392E9, 1.66894644E9, 1.668946488E9, 1.668946536E9, 1.668946584E9, 1.668946632E9, 1.66894668E9, 1.668946728E9, 1.668946776E9, 1.668946824E9, 1.668946872E9, 1.66894692E9, 1.668946968E9, 1.668947016E9, 1.668947064E9, 1.668947112E9, 1.66894716E9, 1.668947208E9, 1.668947256E9, 1.668947304E9, 1.668947352E9, 1.6689474E9, 1.668947448E9, 1.668947496E9, 1.668947544E9, 1.668947592E9, 1.66894764E9, 1.66894794E9, 1.66894812E9, 1.668953962E9, 1.66895401E9, 1.668954058E9, 1.668954106E9, 1.668954154E9, 1.668954202E9, 1.66895425E9, 1.668954298E9, 1.668954346E9, 1.668954394E9, 1.668954442E9, 1.66895449E9, 1.668954538E9, 1.668954586E9, 1.668954634E9, 1.668954682E9, 1.66895473E9, 1.668954778E9, 1.668954826E9, 1.668954874E9, 1.668954922E9, 1.66895497E9, 1.668955018E9, 1.668955066E9, 1.668955114E9, 1.668955162E9, 1.66895521E9, 1.668955258E9, 1.668955306E9, 1.668955354E9, 1.668955402E9, 1.66895545E9, 1.668955498E9, 1.668955546E9, 1.668955594E9, 1.668955642E9, 1.66895569E9, 1.668955738E9, 1.668955786E9, 1.668955834E9, 1.668955882E9, 1.66895593E9, 1.668955978E9, 1.668956026E9, 1.668956074E9, 1.668956122E9, 1.66895617E9, 1.668956218E9, 1.668956266E9, 1.668956314E9, 1.668956362E9, 1.66895641E9, 1.668956458E9, 1.668956506E9, 1.668956554E9, 1.668956602E9, 1.66895665E9, 1.668956698E9, 1.668956746E9, 1.668956794E9, 1.668956842E9, 1.66895689E9, 1.668956938E9, 1.668956986E9, 1.668957034E9, 1.668957082E9, 1.66895713E9, 1.668957178E9, 1.668957226E9, 1.668957274E9, 1.668957322E9, 1.66895737E9, 1.668957418E9, 1.668957466E9, 1.668957514E9, 1.668957562E9, 1.66895761E9, 1.6689579E9, 1.66895808E9, 1.668964026E9, 1.668964074E9, 1.668964122E9, 1.66896417E9, 1.668964218E9, 1.668964266E9, 1.668964314E9, 1.668964362E9, 1.66896441E9, 1.668964458E9, 1.668964506E9, 1.668964554E9, 1.668964602E9, 1.66896465E9, 1.668964698E9, 1.668964746E9, 1.668964794E9, 1.668964842E9, 1.66896489E9, 1.668964938E9, 1.668964986E9, 1.668965034E9, 1.668965082E9, 1.66896513E9, 1.668965178E9, 1.668965226E9, 1.668965274E9, 1.668965322E9, 1.66896537E9, 1.668965418E9, 1.668965466E9, 1.668965514E9, 1.668965562E9, 1.66896561E9, 1.668965658E9, 1.668965706E9, 1.668965754E9, 1.668965802E9, 1.66896585E9, 1.668965898E9, 1.668965946E9, 1.668965994E9, 1.668966042E9, 1.66896609E9, 1.668966138E9, 1.668966186E9, 1.668966234E9, 1.668966282E9, 1.66896633E9, 1.668966378E9, 1.668966426E9, 1.668966474E9, 1.668966522E9, 1.66896657E9, 1.668966618E9, 1.668966666E9, 1.668966714E9, 1.668966762E9, 1.66896681E9, 1.668966858E9, 1.668966906E9, 1.668966954E9, 1.668967002E9, 1.66896705E9, 1.668967098E9, 1.668967146E9, 1.668967194E9, 1.668967242E9, 1.66896729E9, 1.668967338E9, 1.668967386E9, 1.668967434E9, 1.668967482E9, 1.66896753E9, 1.6689678E9, 1.66896798E9, 1.668973745E9, 1.668973793E9, 1.668973841E9, 1.668973889E9, 1.668973937E9, 1.668973985E9, 1.668974033E9, 1.668974081E9, 1.668974129E9, 1.668974177E9, 1.668974225E9, 1.668974273E9, 1.668974321E9, 1.668974369E9, 1.668974417E9, 1.668974465E9, 1.668974513E9, 1.668974561E9, 1.668974609E9, 1.668974657E9, 1.668974705E9, 1.668974753E9, 1.668974801E9, 1.668974849E9, 1.668974897E9, 1.668974945E9, 1.668974993E9, 1.668975041E9, 1.668975089E9, 1.668975137E9, 1.668975185E9, 1.668975233E9, 1.668975281E9, 1.668975329E9, 1.668975377E9, 1.668975425E9, 1.668975473E9, 1.668975521E9, 1.668975569E9, 1.668975617E9, 1.668975665E9, 1.668975713E9, 1.668975761E9, 1.668975809E9, 1.668975857E9, 1.668975905E9, 1.668975953E9, 1.668976001E9, 1.668976049E9, 1.668976097E9, 1.668976145E9, 1.668976193E9, 1.668976241E9, 1.668976289E9, 1.668976337E9, 1.668976385E9, 1.668976433E9, 1.668976481E9, 1.668976529E9, 1.668976577E9, 1.668976625E9, 1.668976673E9, 1.668976721E9, 1.668976769E9, 1.668976817E9, 1.668976865E9, 1.668976913E9, 1.668976961E9, 1.668977009E9, 1.668977057E9, 1.668977105E9, 1.668977153E9, 1.668977201E9, 1.668977249E9, 1.66897752E9, 1.6689777E9, 1.668983522E9, 1.66898357E9, 1.668983618E9, 1.668983666E9, 1.668983714E9, 1.668983762E9, 1.66898381E9, 1.668983858E9, 1.668983906E9, 1.668983954E9, 1.668984002E9, 1.66898405E9, 1.668984098E9, 1.668984146E9, 1.668984194E9, 1.668984242E9, 1.66898429E9, 1.668984338E9, 1.668984386E9, 1.668984434E9, 1.668984482E9, 1.66898453E9, 1.668984578E9, 1.668984626E9, 1.668984674E9, 1.668984722E9, 1.66898477E9, 1.668984818E9, 1.668984866E9, 1.668984914E9, 1.668984962E9, 1.66898501E9, 1.668985058E9, 1.668985106E9, 1.668985154E9, 1.668985202E9, 1.66898525E9, 1.668985298E9, 1.668985346E9, 1.668985394E9, 1.668985442E9, 1.66898549E9, 1.668985538E9, 1.668985586E9, 1.668985634E9, 1.668985682E9, 1.66898573E9, 1.668985778E9, 1.668985826E9, 1.668985874E9, 1.668985922E9, 1.66898597E9, 1.668986018E9, 1.668986066E9, 1.668986114E9, 1.668986162E9, 1.66898621E9, 1.668986258E9, 1.668986306E9, 1.668986354E9, 1.668986402E9, 1.66898645E9, 1.668986498E9, 1.668986546E9, 1.668986594E9, 1.668986642E9, 1.66898669E9, 1.668986738E9, 1.668986786E9, 1.668986834E9, 1.668986882E9, 1.66898693E9, 1.668986978E9, 1.668987026E9, 1.668987074E9, 1.668987122E9, 1.66898717E9, 1.66898742E9, 1.66898772E9, 1.668993676E9, 1.668993724E9, 1.668993772E9, 1.66899382E9, 1.668993868E9, 1.668993916E9, 1.668993964E9, 1.668994012E9, 1.66899406E9, 1.668994108E9, 1.668994156E9, 1.668994204E9, 1.668994252E9, 1.6689943E9, 1.668994348E9, 1.668994396E9, 1.668994444E9, 1.668994492E9, 1.66899454E9, 1.668994588E9, 1.668994636E9, 1.668994684E9, 1.668994732E9, 1.66899478E9, 1.668994828E9, 1.668994876E9, 1.668994924E9, 1.668994972E9, 1.66899502E9, 1.668995068E9, 1.668995116E9, 1.668995164E9, 1.668995212E9, 1.66899526E9, 1.668995308E9, 1.668995356E9, 1.668995404E9, 1.668995452E9, 1.6689955E9, 1.668995548E9, 1.668995596E9, 1.668995644E9, 1.668995692E9, 1.66899574E9, 1.668995788E9, 1.668995836E9, 1.668995884E9, 1.668995932E9, 1.66899598E9, 1.668996028E9, 1.668996076E9, 1.668996124E9, 1.668996172E9, 1.66899622E9, 1.668996268E9, 1.668996316E9, 1.668996364E9, 1.668996412E9, 1.66899646E9, 1.668996508E9, 1.668996556E9, 1.668996604E9, 1.668996652E9, 1.6689967E9, 1.668996748E9, 1.668996796E9, 1.668996844E9, 1.668996892E9, 1.66899694E9, 1.668996988E9, 1.668997036E9, 1.668997084E9, 1.668997132E9, 1.66899718E9, 1.6689975E9, 1.66899768E9, 1.669003569E9, 1.669003617E9, 1.669003665E9, 1.669003713E9, 1.669003761E9, 1.669003809E9, 1.669003857E9, 1.669003905E9, 1.669003953E9, 1.669004001E9, 1.669004049E9, 1.669004097E9, 1.669004145E9, 1.669004193E9, 1.669004241E9, 1.669004289E9, 1.669004337E9, 1.669004385E9, 1.669004433E9, 1.669004481E9, 1.669004529E9, 1.669004577E9, 1.669004625E9, 1.669004673E9, 1.669004721E9, 1.669004769E9, 1.669004817E9, 1.669004865E9, 1.669004913E9, 1.669004961E9, 1.669005009E9, 1.669005057E9, 1.669005105E9, 1.669005153E9, 1.669005201E9, 1.669005249E9, 1.669005297E9, 1.669005345E9, 1.669005393E9, 1.669005441E9, 1.669005489E9, 1.669005537E9, 1.669005585E9, 1.669005633E9, 1.669005681E9, 1.669005729E9, 1.669005777E9, 1.669005825E9, 1.669005873E9, 1.669005921E9, 1.669005969E9, 1.669006017E9, 1.669006065E9, 1.669006113E9, 1.669006161E9, 1.669006209E9, 1.669006257E9, 1.669006305E9, 1.669006353E9, 1.669006401E9, 1.669006449E9, 1.669006497E9, 1.669006545E9, 1.669006593E9, 1.669006641E9, 1.669006689E9, 1.669006737E9, 1.669006785E9, 1.669006833E9, 1.669006881E9, 1.669006929E9, 1.66900722E9, 1.6690074E9, 1.669013278E9, 1.669013326E9, 1.669013374E9, 1.669013422E9, 1.66901347E9, 1.669013518E9, 1.669013566E9, 1.669013614E9, 1.669013662E9, 1.66901371E9, 1.669013758E9, 1.669013806E9, 1.669013854E9, 1.669013902E9, 1.66901395E9, 1.669013998E9, 1.669014046E9, 1.669014094E9, 1.669014142E9, 1.66901419E9, 1.669014238E9, 1.669014286E9, 1.669014334E9, 1.669014382E9, 1.66901443E9, 1.669014478E9, 1.669014526E9, 1.669014574E9, 1.669014622E9, 1.66901467E9, 1.669014718E9, 1.669014766E9, 1.669014814E9, 1.669014862E9, 1.66901491E9, 1.669014958E9, 1.669015006E9, 1.669015054E9, 1.669015102E9, 1.66901515E9, 1.669015198E9, 1.669015246E9, 1.669015294E9, 1.669015342E9, 1.66901539E9, 1.669015438E9, 1.669015486E9, 1.669015534E9, 1.669015582E9, 1.66901563E9, 1.669015678E9, 1.669015726E9, 1.669015774E9, 1.669015822E9, 1.66901587E9, 1.669015918E9, 1.669015966E9, 1.669016014E9, 1.669016062E9, 1.66901611E9, 1.669016158E9, 1.669016206E9, 1.669016254E9, 1.669016302E9, 1.66901635E9, 1.669016398E9, 1.669016446E9, 1.669016494E9, 1.669016542E9, 1.66901659E9, 1.669016638E9, 1.669016686E9, 1.669016734E9, 1.669016782E9, 1.66901683E9, 1.66901724E9, 1.66901742E9, 1.669023366E9, 1.669023414E9, 1.669023462E9, 1.66902351E9, 1.669023558E9, 1.669023606E9, 1.669023654E9, 1.669023702E9, 1.66902375E9, 1.669023798E9, 1.669023846E9, 1.669023894E9, 1.669023942E9, 1.66902399E9, 1.669024038E9, 1.669024086E9, 1.669024134E9, 1.669024182E9, 1.66902423E9, 1.669024278E9, 1.669024326E9, 1.669024374E9, 1.669024422E9, 1.66902447E9, 1.669024518E9, 1.669024566E9, 1.669024614E9, 1.669024662E9, 1.66902471E9, 1.669024758E9, 1.669024806E9, 1.669024854E9, 1.669024902E9, 1.66902495E9, 1.669024998E9, 1.669025046E9, 1.669025094E9, 1.669025142E9, 1.66902519E9, 1.669025238E9, 1.669025286E9, 1.669025334E9, 1.669025382E9, 1.66902543E9, 1.669025478E9, 1.669025526E9, 1.669025574E9, 1.669025622E9, 1.66902567E9, 1.669025718E9, 1.669025766E9, 1.669025814E9, 1.669025862E9, 1.66902591E9, 1.669025958E9, 1.669026006E9, 1.669026054E9, 1.669026102E9, 1.66902615E9, 1.669026198E9, 1.669026246E9, 1.669026294E9, 1.669026342E9, 1.66902639E9, 1.669026438E9, 1.669026486E9, 1.669026534E9, 1.669026582E9, 1.66902663E9, 1.669026678E9, 1.669026726E9, 1.669026774E9, 1.669026822E9, 1.66902687E9, 1.6690272E9}
    LATITUDE = 
      {38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2545, 38.2572, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.257, 38.26, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2637, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2638, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2635, 38.2632, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.263, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2627, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2615, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.2612, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.261, 38.2603, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2588, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2585, 38.2592, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2587, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2602, 38.2605, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.26, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.2598, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.259, 38.2568, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2565, 38.2525, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.2507, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.243, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2433, 38.2663, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2665, 38.2877, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.2878, 38.3088, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.309, 38.3295, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3298, 38.3493, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.349, 38.3583, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3578, 38.3678, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3673, 38.3752, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.375, 38.38, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3798, 38.3843, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3842, 38.3887, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3885, 38.3927, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3955, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.3953, 38.399, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.3985, 38.4015, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4012, 38.4047, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4043, 38.4073, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.407, 38.4105, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4102, 38.4128, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4127, 38.4145, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.414, 38.4173, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4168, 38.4205, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.423, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4225, 38.4253, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4248, 38.4272, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4267, 38.4295, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.429, 38.4322, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4317, 38.4357, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4353, 38.4382, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4413, 38.4463, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4467, 38.4507, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4508, 38.4535, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4537, 38.4562, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4563, 38.4593, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4597, 38.4632, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4635, 38.4672, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4673, 38.4705, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.471, 38.4745, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4748, 38.4783, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4787, 38.4817, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.4822, 38.485, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4853, 38.4877, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.488, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.4895, 38.491, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.4912, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.492311111111114, 38.4932, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.493, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.494238461538465, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.4953, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.49685769230769, 38.498, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.4978, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.499144, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.49825, 38.4963, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.4965, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.49432222222222, 38.4923, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.4925, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.48972222222222, 38.4875, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.4877, 38.485, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4852, 38.4823, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4827, 38.4802, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4803, 38.4768, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.477, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4738, 38.4702, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.47, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4668, 38.4632, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4633, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.4605, 38.458, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4582, 38.4553, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4555, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4528, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4503, 38.4473, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4472, 38.4442, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.444, 38.441, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4407, 38.4382, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.4378, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.435, 38.4317, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4312, 38.4275, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4268, 38.4242, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4238, 38.4212, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4207, 38.4172, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4167, 38.4127, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.412, 38.4083, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4078, 38.4043, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.404, 38.3983, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.3978, 38.392, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3915, 38.3832, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3828, 38.3722, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.372, 38.36, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3597, 38.3492, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3487, 38.3337, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3333, 38.3158, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.315, 38.2988, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.298, 38.285, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2842, 38.2693, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2687, 38.2533, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.24, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2393, 38.2297, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.229, 38.2183, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2178, 38.2053, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.2047, 38.1923, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1917, 38.1812, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1807, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1712, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1578, 38.1458, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1455, 38.1363, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1362, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1315, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.1205, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.094, 38.0855, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0852, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0747, 38.0622, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0618, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.0488, 38.039, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0392, 38.0308, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.031, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0178, 38.0003, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9998, 37.9862, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.9858, 37.976, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.9758, 37.965, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9652, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9498, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9327, 37.9193, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.919, 37.9088, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.9087, 37.8937, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8932, 37.8745, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8742, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8557, 37.8408, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.84, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.827, 37.8105, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.8103, 37.7897, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7895, 37.7698, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7697, 37.7562, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7558, 37.7403, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7398, 37.7173, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.7168, 37.6942, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6937, 37.6787, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.678, 37.6657, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6652, 37.6482, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6478, 37.6265, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6257, 37.6067, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.606, 37.5907, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5902, 37.5762, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5758, 37.5558, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.5553, 37.531, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5308, 37.5058, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.5055, 37.4845, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4842, 37.4657, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4655, 37.4492, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.449, 37.4298, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4292, 37.4143, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4142, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.4032, 37.3948, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.395, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3867, 37.3778, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.378, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3692, 37.3627, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.363, 37.355, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3558, 37.3522, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.3527, 37.345, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3457, 37.3412, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3418, 37.3362, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3365, 37.3263, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3265, 37.3123, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3127, 37.3003, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.3007, 37.2903, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2908, 37.2792, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.2795, 37.268, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2683, 37.2568, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2572, 37.2448, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2452, 37.2558, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2563, 37.2658, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.266, 37.2782, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2783, 37.2912, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.2915, 37.3105, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.3108, 37.331, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3312, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3483, 37.3673, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3678, 37.3923, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.3927, 37.4162, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4383, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4525, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4762, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.4847, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.488, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.49, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4948, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4987, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.5023, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.4985, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.493, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4888, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.4918, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4958, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.496, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4992, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.5035, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.509, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5093, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.508, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5087, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.524, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5267, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.5288, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5348, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5515, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.5593, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5635, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.584, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6417, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.661, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.673, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6923, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.7083, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7202, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7317, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7455, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7852, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.798, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.8133, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8273, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8373, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.8443, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.857, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8728, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8862, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.8948, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9503, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9695, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9693, 37.9828, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9825, 37.9978, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 37.998, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0098, 38.0208, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.021, 38.0347, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0348, 38.0533, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0535, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0703, 38.0813, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0812, 38.0983, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.0987, 38.1167, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.117, 38.1378, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.138, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.156, 38.1732, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.173, 38.191, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.1907, 38.2105, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2107, 38.2342, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2347, 38.2522, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.2527, 38.262, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.2623, 38.276, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2762, 38.2958, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.2957, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3145, 38.3273, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.327, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3387, 38.3558, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3555, 38.3713, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3708, 38.3808, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.3807, 38.386, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3857, 38.3877, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3878, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3873, 38.3885, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3877, 38.3898, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3892, 38.3912, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.3905, 38.392, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3913, 38.3937, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.3928, 38.395, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3952, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3943, 38.3953, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3953, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3947, 38.3965, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3958, 38.3977, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.397, 38.3988, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.3982, 38.4005, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.3997, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.401900000000005, 38.404, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.404336585365854, 38.4058, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4073, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.4063, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.407560000000004, 38.4087, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.4073, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.407250000000005, 38.4072, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.4057, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.40595641025641, 38.4062, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.4052, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40553333333333, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.40586666666667, 38.4062, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.4055, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.40752692307693, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.409792307692314, 38.4117, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.4112, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41207962962963, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.41295925925926, 38.4137, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.4132, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.41752777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.42162777777778, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.4255, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.42958, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.43366, 38.4375, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.437, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44092727272727, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.44460909090909, 38.4478, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.4473, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.45144375, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.4555875, 38.459, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.4588, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46236666666666, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.46617111111111, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.4695, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.47340697674418, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.476825581395346, 38.48, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.4805, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.48378666666667, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.486686666666664, 38.4892, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.4898, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49163333333333, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.49359761904762, 38.4953, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.4955, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.496433333333336, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.49751025641026, 38.4983, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.4987, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.49911219512195, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.499524390243906, 38.5, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.5002, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.498066666666666, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.495780952380954, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4938, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4907, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4876, 38.4845, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.4848, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.480533333333334, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.47626666666667, 38.472, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4722, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.4671, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.462, 38.4572, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.457, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.45243076923077, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.44786153846154, 38.4438, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.4435, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43933965517241, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.43517931034483, 38.4308, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.4298, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.42518, 38.421, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.4202, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.41534893617021, 38.4107, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.41, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.40665, 38.4033, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.4028, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.40075, 38.3987, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.396058823529415, 38.394, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.3937, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.39326607142857, 38.3928, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.3923, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.389989743589744, 38.387, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3868, 38.3778, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3777, 38.3657, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3655, 38.3563, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.3565, 38.348, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3482, 38.3407, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.341, 38.3335, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3338, 38.3248, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3252, 38.3137, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3138, 38.3062, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3057, 38.3012, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.3013, 38.2987, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.299, 38.293, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2933, 38.2837, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.2838, 38.28, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2803, 38.2762, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2765, 38.2703, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2708, 38.2625, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2628, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2557, 38.2527, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.2488, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.2445, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.242, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2427, 38.2383, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2388, 38.2348, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2355, 38.2303, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2308, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2215, 38.2133, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2135, 38.2072, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2073, 38.2017, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.2015, 38.1962, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.196, 38.1923, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1927, 38.1897, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1902, 38.1853, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1857, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1795, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1723, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.1673, 38.162, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1618, 38.1548, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.1543, 38.15, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1493, 38.1458, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1457, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1427, 38.1365, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1358, 38.1322, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1317, 38.1078, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.107, 38.0812, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0808, 38.0545, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.0543, 38.04, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0398, 38.0273, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.0268, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.016, 38.0043, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 38.0038, 37.9985, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9983, 37.9923, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.9925, 37.988, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9882, 37.9808, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9805, 37.9722, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.9717, 37.965, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.9645, 37.961, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.9607, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.956, 37.9488, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9485, 37.9403, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9398, 37.9342, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9338, 37.9295, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.9293, 37.923, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9228, 37.9132, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.913, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.906, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.9005, 37.8957, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8958, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.8875, 37.876, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8758, 37.8683, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8682, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.8647, 37.858, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.8578, 37.847, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8468, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8355, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8317, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.8273, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.816, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.8048, 37.795, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7955, 37.7895, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.7897, 37.781, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7807, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.7693, 37.761}
    LONGITUDE = 
      {-123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.3333, -123.337, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3417, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3415, -123.3473, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3472, -123.3547, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.361, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3608, -123.3685, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.3682, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.376, -123.384, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3837, -123.3907, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.39, -123.3953, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.3947, -123.4, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.3995, -123.4062, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4138, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4135, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4235, -123.4367, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.437, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4528, -123.4693, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4692, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.4862, -123.5075, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.5077, -123.533, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5332, -123.5593, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5602, -123.5688, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.569, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.58, -123.591, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.5907, -123.6012, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.6008, -123.613, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.6135, -123.5942, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5948, -123.5777, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.5778, -123.565, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5652, -123.5545, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5547, -123.5457, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.546, -123.537, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5372, -123.5283, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5285, -123.5202, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.5207, -123.513, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.5135, -123.508, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5083, -123.5018, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.5022, -123.4958, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.496, -123.4888, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.489, -123.4817, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.4813, -123.473, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4723, -123.4665, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4662, -123.4612, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.4552, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.455, -123.4495, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4493, -123.4442, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4443, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4398, -123.4352, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4353, -123.4305, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4308, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.422, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4222, -123.4157, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.416, -123.41, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4103, -123.4053, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4022, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.4025, -123.3977, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.398, -123.3932, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3935, -123.3893, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.3898, -123.386, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3863, -123.3827, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3828, -123.3787, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3788, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3742, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.365, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3648, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3605, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.3562, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35275555555555, -123.35, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.3502, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.34696923076923, -123.3442, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.3443, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.34164615384616, -123.3397, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.3402, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.338016, -123.3363, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3368, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.3434, -123.35, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.3505, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.35775925925927, -123.3645, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.365, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.37238888888888, -123.3783, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3787, -123.3852, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3857, -123.3907, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3903, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3942, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.3993, -123.4055, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4058, -123.4123, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4125, -123.4193, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4197, -123.4263, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4262, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4323, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.4383, -123.444, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4435, -123.4492, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.449, -123.4557, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.462, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4618, -123.4682, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4678, -123.4743, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4815, -123.4882, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4877, -123.4928, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4925, -123.4987, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.4982, -123.5057, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5053, -123.5133, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5128, -123.5212, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5205, -123.5287, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5282, -123.5378, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5377, -123.5478, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5475, -123.5572, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.557, -123.5677, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.5675, -123.583, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.5828, -123.6022, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.602, -123.629, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6288, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6617, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.6922, -123.7208, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7207, -123.7517, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7518, -123.7842, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.7847, -123.8162, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.8163, -123.846, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8462, -123.8742, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.8743, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.902, -123.9313, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.9315, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.962, -123.9895, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -124.0178, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.018, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0472, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.0753, -124.1018, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1022, -124.1297, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.1302, -124.159, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1597, -124.1862, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.1868, -124.2122, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2127, -124.2378, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2382, -124.2642, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2645, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.2942, -124.3228, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3238, -124.3533, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.354, -124.3825, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.383, -124.4102, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.4108, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.435, -124.4603, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4605, -124.4918, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.4927, -124.5263, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5273, -124.5592, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5598, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.5872, -124.614, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6142, -124.6457, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.6462, -124.682, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.6825, -124.7168, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.7173, -124.75, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7503, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.8233, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8243, -124.8613, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8622, -124.8967, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.8972, -124.9297, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.93, -124.9663, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -124.9665, -125.006, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.0062, -125.042, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0423, -125.0763, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.0767, -125.1138, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1143, -125.1537, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.154, -125.19, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.1905, -125.2265, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2272, -125.2638, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.2645, -125.3007, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.3012, -125.337, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3373, -125.3728, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.3732, -125.4077, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.408, -125.4413, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4417, -125.4752, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.4755, -125.5138, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.5143, -125.564, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.5645, -125.6193, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6198, -125.6707, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.6712, -125.7228, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7233, -125.7787, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.7793, -125.8322, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.833, -125.8737, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.8742, -125.9073, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9078, -125.9417, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9423, -125.9805, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -125.9817, -126.0152, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.0163, -126.043, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0437, -126.0672, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.068, -126.0957, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.0968, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1158, -126.1275, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1278, -126.1375, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.138, -126.1462, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1467, -126.1588, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.1592, -126.167, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1672, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1712, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1718, -126.1802, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1798, -126.1558, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1555, -126.1345, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1343, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.1113, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0897, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0752, -126.0575, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0573, -126.0395, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0393, -126.0225, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.023, -126.0132, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0133, -126.0027, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9623, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9347, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9088, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.8858, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8582, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8303, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8092, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.7898, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.774, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7555, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7413, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7318, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7292, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7232, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7083, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.6978, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6907, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.6828, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.67, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6578, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6512, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6473, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6337, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6187, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6025, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.5942, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.569, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.4938, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.425, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.3993, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3705, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3012, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.2605, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.2253, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1592, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.0763, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0393, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0087, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -124.976, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9457, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.915, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.8817, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.846, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8135, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.7847, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7602, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7333, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.6717, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.64, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.609, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.5815, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5177, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4875, -124.4557, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.456, -124.4285, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4288, -124.4005, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.4007, -124.3677, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3675, -124.3312, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.3308, -124.2968, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.2965, -124.258, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2575, -124.2218, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.2213, -124.188, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1875, -124.1468, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.1458, -124.107, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.106, -124.066, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0263, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -124.0253, -123.9905, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9898, -123.9548, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.9542, -123.918, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.9177, -123.8787, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.878, -123.837, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.836, -123.7975, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7967, -123.7625, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.7272, -123.6947, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6943, -123.6627, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.662, -123.6308, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.63, -123.6033, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.6027, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5843, -123.5712, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5708, -123.5602, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5595, -123.5487, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.548, -123.5395, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.539, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5333, -123.5278, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5277, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5228, -123.5203, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5208, -123.5183, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5188, -123.5173, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5178, -123.5163, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5165, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.5137, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.511, -123.5067, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5065, -123.5012, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.5007, -123.4957, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.4953, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.49064418604651, -123.4862, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.4857, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.48267804878049, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.4798, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.47754761904761, -123.4755, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4757, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4736, -123.4717, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.472, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.469, -123.466, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.4665, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.46342307692308, -123.4605, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.461, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45706666666666, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.45313333333334, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.4492, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44629038461538, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.44303846153846, -123.4403, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.4405, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.43476481481481, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.42902962962962, -123.4242, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.4245, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.42126296296296, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4181962962963, -123.4153, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.4148, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.41021, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.40562, -123.4013, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.4007, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39608181818183, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.39175227272727, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.388, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38552083333333, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.38304166666667, -123.381, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.3815, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37966666666667, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.37771111111111, -123.376, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.3768, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37508837209303, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.37359069767443, -123.3722, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.3733, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37216666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.37116666666667, -123.3703, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3708, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.3698, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.36872857142858, -123.3678, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.3688, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36793333333333, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.36693333333334, -123.3662, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.3672, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.36643902439025, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3656780487805, -123.3648, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.3653, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37193333333333, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.37904047619048, -123.3852, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.386, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39266666666667, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.39933333333333, -123.406, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.4073, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41363333333334, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.41996666666667, -123.4263, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.4265, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.433402, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.440304, -123.4468, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.447, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.45433846153846, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.46167692307692, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.4682, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.47478448275862, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.48136896551723, -123.4883, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.487, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4914625, -123.4955, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.4943, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.49940638297872, -123.5043, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.5035, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.51085, -123.5182, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.5175, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.52525, -123.533, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.53903921568627, -123.546, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.545, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.55319642857143, -123.562, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.5613, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.57394102564103, -123.5903, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.5897, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6042, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.6212, -123.644, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.6442, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.666, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.6867, -123.7025, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7022, -123.7155, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7148, -123.7295, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7287, -123.7457, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.745, -123.7622, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7617, -123.7798, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7797, -123.7943, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.7945, -123.8078, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8072, -123.8232, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8227, -123.8347, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.834, -123.8452, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.845, -123.8532, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.852, -123.8642, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8632, -123.8733, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.873, -123.8833, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.882, -123.8915, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.8907, -123.9057, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.9052, -123.915, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.9137, -123.917, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9162, -123.9253, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.925, -123.9393, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.939, -123.9532, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9527, -123.9638, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.963, -123.9713, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9702, -123.9818, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.981, -123.9973, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -123.9968, -124.0115, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0105, -124.0163, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.015, -124.0257, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.025, -124.0388, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0383, -124.0543, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0537, -124.0655, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0647, -124.0725, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.0715, -124.079, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0778, -124.0922, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.0917, -124.1065, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.1057, -124.115, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1138, -124.1218, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.121, -124.1178, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1165, -124.1142, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1133, -124.1107, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1098, -124.1187, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.118, -124.1303, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1298, -124.1435, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1432, -124.1568, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1563, -124.1713, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.171, -124.1883, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.188, -124.208, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2077, -124.2275, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.227, -124.2433, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2428, -124.2587, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2583, -124.2743, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.274, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.2938, -124.315, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3147, -124.3375, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.3373, -124.358, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3578, -124.3785, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3783, -124.3985, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.3982, -124.4187, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.4182, -124.439, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.4387, -124.458, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4577, -124.4782, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4778, -124.4985, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.4982, -124.5197, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.5195, -124.541, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5407, -124.5622, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5618, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.5843, -124.6035, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6033, -124.6275, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.6277, -124.657, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6572, -124.6828, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.6827, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.7042, -124.729, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7292, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.7558, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.78, -124.804, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8042, -124.8302, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8303, -124.8602}
    DEPTH = 
      {NaN, 105.732895, 105.336105, 104.780594, 104.10604, 103.31245, 102.598206, 101.84429, 100.85229, 100.13804, 98.86826, 98.233376, 96.884224, 95.733475, 94.74144, 93.511314, 92.24149, 89.90025, 88.74946, 86.328804, 84.979576, 83.51129, 82.12236, 80.85248, 79.344475, 77.4793, 76.24907, 74.50292, 73.312355, 72.00273, 70.335915, 69.065956, 67.59756, 65.77196, 64.46229, 62.795414, 61.565094, 60.096638, 58.509106, 57.239075, 55.810276, 54.024265, 52.635136, 50.92848, 49.658394, 48.189854, 46.52285, 45.17336, 43.74448, 42.11713, 40.886684, 39.25931, 38.028854, 36.599922, 34.853436, 33.662643, 32.23368, 30.72532, 29.494808, 28.1849, 26.676512, 25.48567, 24.175735, 22.667316, 21.198584, 20.166492, 18.69774, 17.467155, 16.157171, 14.648693, 13.497479, 12.227166, 10.718659, 9.567423, 7.9795, 6.3915644, 5.319701, 3.771444, 2.54077, 1.4688865, NaN, NaN, 108.5104, 108.23265, 107.67715, 107.08196, 106.2487, 105.45512, 104.74088, 103.59018, 102.875946, 101.80458, 100.852264, 99.89993, 98.9476, 98.03494, 97.0826, 96.050896, 94.423965, 93.07479, 91.36847, 90.09864, 88.63039, 87.32086, 86.051, 84.543045, 82.51918, 81.16993, 79.66193, 77.87613, 76.48716, 74.7807, 73.471085, 72.0424, 69.97872, 68.669075, 66.88318, 65.6132, 64.10509, 62.319145, 60.96976, 59.223484, 57.83439, 56.365906, 54.381454, 53.270153, 51.52381, 50.214046, 48.7852, 47.15789, 45.808403, 44.538292, 42.791874, 41.521744, 39.735607, 38.386074, 37.15561, 35.40913, 34.09926, 32.868767, 31.161945, 29.931435, 28.581837, 26.835283, 25.604748, 23.93756, 22.66731, 21.476446, 19.84892, 18.618343, 17.228973, 15.7602005, 14.608993, 13.29899, 11.830189, 10.639261, 8.971951, 7.423722, 6.2327685, 4.962411, 3.533249, 2.4216714, 1.15129, NaN, NaN, 126.08729, 124.9367, 123.31, 121.762634, 120.33429, 118.310776, 116.247574, 114.10499, 110.930756, 107.558075, 104.82021, 102.08231, 98.66981, 95.53501, 92.51922, 89.46369, 86.40813, 83.43188, 80.45559, 77.3602, 74.38382, 71.44709, 68.47062, 65.49412, 62.75569, 59.818787, 57.159664, 54.659264, 51.920692, 49.102707, 46.36406, 43.34754, 40.291283, 37.6716, 34.972496, 32.074886, 29.296322, 26.597107, 23.858162, 21.11918, 18.340466, 15.482319, 12.703527, 10.162885, 7.1855297, 4.4066253, 1.9055793, NaN, NaN, 131.60207, 130.4912, 129.18193, 127.59493, 125.8889, 124.18285, 122.19906, 120.05654, 117.08078, 113.86691, 111.32753, 108.78811, 105.65347, 102.99494, 100.17766, 97.24129, 94.066795, 90.89225, 88.0748, 85.29699, 82.55883, 79.78095, 77.16177, 74.30444, 71.685196, 69.14529, 66.406906, 63.708183, 61.168175, 58.310627, 55.611794, 52.952618, 49.737743, 47.15787, 44.260437, 40.96604, 37.55252, 34.41679, 31.638256, 28.81999, 25.763517, 23.143646, 20.404655, 17.864109, 15.32353, 12.822618, 10.162884, 7.344322, 4.92271, 2.3819714, NaN, NaN, 134.29991, 133.26839, 131.87979, 130.37218, 128.82486, 127.07916, 125.17475, 123.19096, 120.175575, 116.76337, 113.90659, 111.208496, 107.63743, 104.344055, 101.52679, 98.43172, 95.41596, 92.36049, 89.38432, 86.56686, 83.94776, 81.20958, 78.630104, 76.01091, 73.27263, 70.69305, 68.11344, 65.25599, 62.239746, 59.66003, 56.961216, 54.460815, 51.92069, 49.142395, 46.324368, 43.585686, 40.45005, 37.631905, 35.012188, 32.511517, 29.891731, 27.271914, 24.81084, 22.230654, 19.848913, 17.268663, 14.886866, 12.4653425, 9.68651, 7.026736, 4.6845174, 2.1834748, NaN, NaN, 138.66397, 137.63248, 136.24391, 134.73633, 133.07002, 131.24501, 129.41998, 127.43624, 124.460594, 121.68328, 119.263016, 116.723694, 114.06531, 111.32754, 108.27229, 105.45508, 102.79655, 100.098305, 97.241295, 94.58266, 91.92399, 89.10655, 86.32876, 83.590614, 80.733376, 77.91579, 75.09815, 72.39954, 69.66121, 66.922844, 64.18444, 61.52537, 58.985332, 56.524643, 53.7861, 51.245964, 48.66611, 45.88777, 43.38723, 40.767586, 37.830368, 35.369423, 32.948143, 30.407753, 27.86733, 25.485655, 23.024563, 20.56344, 17.983198, 15.402925, 12.981408, 10.361374, 7.622211, 5.2403007, 2.6995654, 1.032191, NaN, NaN, 140.88565, 139.73515, 138.26726, 136.68033, 134.9347, 133.18904, 131.20534, 129.02324, 126.52372, 123.905136, 121.60393, 119.263016, 116.92208, 114.303375, 111.525925, 108.86748, 106.288345, 103.55047, 100.93159, 98.511086, 95.7731, 93.35253, 90.97162, 88.550995, 86.05098, 83.3922, 80.61433, 77.91579, 74.9791, 72.20112, 69.34373, 66.72441, 63.787563, 61.049118, 58.350323, 55.572113, 52.793865, 50.25372, 47.55478, 44.93519, 42.315563, 39.537136, 36.560207, 33.821396, 31.082548, 28.264273, 25.68413, 23.22304, 20.523745, 18.062592, 15.601409, 12.981408, 10.5201645, 6.907641, 4.3669267, 2.0246775, NaN, NaN, 144.69418, 143.58337, 142.23453, 140.72697, 139.06071, 137.19609, 135.45047, 133.2684, 130.25317, 126.84113, 124.18288, 121.3262, 117.71564, 114.739845, 111.80369, 108.867485, 106.12964, 103.27272, 100.49512, 97.638115, 94.5033, 91.606544, 88.67005, 85.85257, 82.83663, 80.098434, 77.36021, 74.820366, 72.32018, 69.74059, 66.92285, 64.303505, 61.803192, 59.02503, 56.44527, 53.825794, 50.888763, 48.11045, 45.53056, 42.95063, 40.053135, 37.393757, 34.81373, 32.114586, 29.534489, 27.113138, 24.572676, 22.190962, 19.690132, 17.189274, 14.847171, 12.346252, 9.32923, 6.4312596, 3.9699373, 1.4291863, NaN, NaN, 150.20848, 149.13737, 147.47119, 146.04303, 144.17845, 142.39322, 140.36993, 138.34662, 135.4108, 132.47493, 129.85643, 127.55529, 124.976395, 122.35779, 119.382065, 116.60468, 113.90662, 111.20852, 108.31199, 105.574135, 102.83624, 100.05864, 97.36035, 94.78108, 91.963684, 89.50339, 86.9637, 84.304924, 81.765175, 79.304756, 76.68557, 74.22509, 71.7249, 68.98656, 66.287865, 63.7082, 60.850685, 58.191574, 55.61181, 52.83356, 50.094967, 47.475407, 44.657356, 42.156803, 39.69591, 37.1556, 34.615265, 31.995506, 29.097855, 26.319248, 23.699385, 20.76192, 18.340467, 15.879288, 13.378382, 10.877445, 8.058892, 5.4784937, 3.3744519, 1.3497874, NaN, NaN, 157.78546, 156.51604, 155.04826, 153.34245, 151.5573, 149.53409, 147.62988, 145.36862, 142.27422, 139.14008, 136.68036, 134.14125, 130.96732, 128.30913, 125.611206, 122.5165, 119.42175, 116.52534, 113.74792, 110.772064, 107.91521, 105.01863, 102.20137, 99.18568, 96.48738, 93.78905, 90.97164, 88.3526, 85.65417, 83.27316, 80.85245, 78.51107, 75.77282, 73.07422, 70.37558, 67.75628, 65.05757, 62.4382, 59.660046, 56.881855, 54.063934, 51.285667, 48.54705, 46.28469, 44.0223, 41.759888, 39.49745, 37.155605, 34.813732, 32.23367, 29.653574, 27.152836, 24.374203, 21.79401, 19.33287, 16.871704, 14.489901, 11.8698845, 8.932252, 5.9151793, 3.5332484, 1.9055798, NaN, NaN, 164.05312, 162.94241, 161.43501, 159.8086, 157.98383, 156.0797, 154.0962, 151.95403, 149.01839, 145.88437, 143.34538, 140.80635, 137.55318, 134.81572, 132.03854, 128.98361, 125.888954, 123.0323, 120.09627, 117.08083, 113.86696, 110.85143, 107.994576, 105.098, 102.122025, 99.185684, 96.32867, 93.35256, 90.21769, 87.36054, 84.46368, 81.76519, 78.82856, 75.891884, 72.99486, 69.7803, 66.76412, 63.7479, 60.96976, 58.032833, 55.214928, 52.476364, 49.658386, 46.602222, 44.220764, 41.601128, 38.94177, 36.441143, 34.09926, 31.598576, 29.058167, 26.319254, 23.540607, 21.0001, 18.340471, 15.720505, 13.378385, 10.917145, 8.297083, 5.954879, 3.4538507, 1.7467823, NaN, NaN, 174.56487, 173.37488, 171.9469, 170.39989, 168.69421, 166.82985, 164.92581, 162.86307, 159.49124, 155.802, 152.98544, 150.20851, 146.75714, 143.50406, 140.4493, 137.15645, 133.86356, 130.80864, 127.55531, 124.341606, 121.36591, 118.39017, 115.216, 111.72436, 109.14526, 106.12966, 103.27274, 100.25706, 97.439735, 94.7811, 91.84466, 89.0669, 86.40816, 83.82874, 81.01119, 78.27297, 75.65378, 72.63769, 69.93904, 67.4388, 64.54165, 61.76352, 58.985355, 56.00871, 52.95264, 50.412495, 47.63418, 44.736748, 42.474342, 39.93407, 37.1953, 34.932816, 32.55122, 30.010824, 27.4307, 24.771156, 22.190968, 19.76953, 17.348063, 14.966266, 12.584439, 10.123191, 7.820705, 5.4784946, 3.1362576, 1.3894871, NaN, NaN, 189.04242, 186.18665, 182.9342, 179.20572, 173.41454, 167.94052, 162.22836, 156.51605, 150.72423, 145.4083, 140.17159, 135.01408, 129.69774, 124.38127, 118.98531, 113.82728, 108.58975, 103.193375, 97.7175, 92.47956, 87.24149, 82.24139, 77.1618, 72.32019, 67.002235, 62.081017, 56.921547, 52.079464, 47.078506, 42.156807, 36.838066, 31.598574, 26.676504, 22.310051, 18.181684, 14.212023, 9.845305, 5.399097, 2.0643773, NaN, NaN, 204.78807, 202.01186, 198.83897, 195.11078, 189.71667, 184.56042, 179.16605, 173.69218, 168.21819, 162.4267, 156.47636, 150.76389, 144.89256, 139.02106, 133.22874, 127.515625, 122.04039, 116.723724, 111.32756, 106.08997, 100.81257, 95.1779, 89.701805, 84.30493, 78.66981, 73.11391, 67.63722, 62.319138, 57.00092, 51.523808, 46.205307, 41.204205, 36.20298, 31.439796, 26.676502, 22.151268, 17.546543, 12.465346, 7.6222124, 2.858363, NaN, NaN, 229.85176, 226.91724, 223.5068, 219.69975, 213.98903, 208.19882, 201.85321, 195.74538, 189.79602, 183.44983, 177.5001, 171.55022, 165.67949, 160.12593, 154.49289, 148.8597, 143.3057, 137.75154, 132.19724, 126.72212, 121.088165, 115.454056, 109.9785, 104.344086, 98.94759, 93.550964, 87.83673, 82.51917, 77.201485, 72.121765, 67.12129, 62.279453, 57.4375, 52.516052, 47.673866, 42.831566, 37.750996, 32.6703, 27.98642, 23.540607, 19.015305, 14.688386, 10.12319, 5.6769876, 2.0643773, NaN, NaN, 262.60443, 259.82898, 256.33978, 252.61264, 247.45796, 242.85829, 237.94128, 232.94485, 227.71037, 222.47575, 217.39963, 212.24406, 207.00905, 201.61526, 196.14201, 190.66861, 185.0364, 179.40405, 174.08887, 168.85287, 163.37875, 157.90448, 151.87468, 146.55878, 141.00471, 136.40265, 131.72115, 127.039536, 122.51652, 117.596634, 112.517914, 107.28036, 101.88394, 96.72548, 91.64625, 86.64625, 81.80487, 77.28085, 72.75674, 68.15315, 63.39071, 58.62816, 53.4686, 48.229534, 43.149097, 37.98915, 33.22601, 28.383366, 23.461218, 18.697737, 13.85475, 8.614668, 3.7714431, 0.83369344, NaN, NaN, 280.64395, 277.86874, 274.37988, 270.49448, 264.54727, 258.75848, 252.65233, 246.78392, 240.59811, 234.41211, 228.30524, 222.03957, 216.01164, 209.98355, 204.35187, 198.40276, 192.77077, 186.74197, 180.6337, 174.44589, 168.33723, 162.06973, 156.27806, 150.56558, 145.01161, 139.06078, 133.34781, 127.79338, 121.921394, 115.89053, 110.0182, 104.5425, 99.22538, 93.67003, 88.11453, 82.32078, 77.08244, 71.84398, 67.00225, 62.160404, 57.120003, 51.960407, 46.880062, 42.037743, 37.036537, 32.03521, 27.271927, 22.349752, 17.348066, 12.505047, 7.582516, 2.898063, NaN, NaN, 307.72015, 305.0246, 301.77402, 297.88913, 292.33914, 287.0269, 281.31802, 275.8469, 270.4549, 264.90417, 259.11542, 253.40579, 247.93391, 242.5412, 236.8311, 231.5174, 226.20357, 221.04822, 215.81343, 210.18192, 204.94684, 199.47368, 193.92104, 188.36824, 182.41867, 176.62756, 170.83632, 165.12422, 159.33264, 153.62024, 148.06636, 142.51233, 137.27554, 132.11797, 126.801544, 121.326294, 115.61283, 109.89921, 104.74094, 99.741264, 94.34465, 89.10663, 84.10657, 79.18576, 74.74105, 70.21688, 65.53386, 60.850727, 56.32625, 51.563526, 47.03884, 42.11714, 37.35409, 32.908478, 28.224602, 23.54062, 19.015314, 14.5693035, 10.202591, 5.676991, 2.5010715, NaN, NaN, 344.5824, 341.9666, 338.79587, 335.14948, 329.9176, 324.76486, 319.29486, 313.9833, 308.83014, 303.35974, 297.73062, 292.10135, 286.31335, 280.76306, 275.4505, 270.45496, 265.22144, 260.14636, 254.75397, 249.20282, 243.61186, 238.13972, 232.58813, 227.03639, 221.72244, 216.48766, 211.25275, 206.09703, 201.0205, 195.70587, 190.54976, 185.47284, 180.23715, 175.2393, 170.08269, 164.92592, 160.00705, 155.24673, 150.40698, 145.5671, 140.6081, 135.68863, 130.68971, 126.00807, 121.16762, 116.247696, 111.32765, 106.32813, 101.24914, 96.328735, 91.32886, 86.32885, 81.32872, 76.64595, 71.64559, 66.9626, 62.51763, 57.993183, 53.6274, 49.42028, 45.014618, 40.251633, 35.60762, 31.320742, 26.954386, 22.508547, 18.419876, 14.291428, 10.004105, 5.915184, 2.501072, NaN, NaN, 399.66528, 397.05017, 393.95956, 390.47263, 385.08365, 379.77377, 373.8297, 368.28177, 362.4959, 356.8684, 351.0822, 345.4544, 340.06424, 334.67395, 329.36276, 324.05145, 318.34363, 312.63562, 306.4518, 300.5056, 294.2025, 288.25598, 282.22998, 276.2831, 270.25677, 264.46817, 258.67938, 253.12834, 247.25993, 241.78789, 236.3157, 230.60544, 224.97432, 219.34306, 214.0289, 208.63528, 202.92426, 197.45103, 191.73969, 186.18683, 180.43552, 174.48569, 168.85304, 163.29958, 157.82529, 152.35086, 146.95563, 141.6396, 136.40279, 131.16583, 126.24615, 121.32635, 116.32707, 111.327675, 106.2488, 101.09044, 95.852585, 90.85269, 85.85267, 80.693794, 75.57448, 70.09785, 64.938576, 59.85855, 54.937157, 50.253784, 45.173393, 40.251644, 35.40916, 31.042892, 26.835308, 22.548246, 18.181704, 13.973854, 9.607127, 5.3197045, 2.3025758, NaN, NaN, 401.64658, 398.95224, 395.70316, 391.58228, 385.79706, 380.56644, 374.7809, 369.233, 363.76422, 358.05746, 352.42984, 346.80206, 341.2534, 335.46677, 329.91782, 324.44797, 318.8194, 313.27, 307.72043, 302.24997, 296.58118, 290.7933, 284.7674, 278.66202, 272.9529, 267.32297, 261.77216, 256.30048, 250.98729, 245.59465, 240.20186, 234.88824, 229.41586, 223.86403, 218.39136, 212.83923, 207.44559, 201.89316, 196.57855, 191.34314, 186.02826, 180.79256, 175.47742, 170.47945, 165.16403, 160.08649, 155.00882, 149.93102, 144.69441, 139.45767, 134.37949, 129.06313, 124.22275, 119.302895, 114.22421, 109.22476, 104.46327, 99.70167, 94.93995, 90.09876, 85.33682, 80.45572, 75.733246, 71.20909, 66.36734, 62.041416, 57.834465, 53.70681, 49.46, 45.2131, 41.204266, 37.076275, 32.9482, 28.82004, 24.929968, 21.000128, 16.911425, 12.902035, 8.138302, 3.8508463, 1.3497895, NaN, NaN, 401.28937, 398.59506, 395.34595, 391.70056, 386.3116, 381.23953, 376.16733, 370.69873, 365.1507, 359.5233, 354.05423, 348.58502, 343.1157, 337.80472, 332.25583, 326.78604, 321.31613, 315.92532, 310.5344, 305.14334, 299.63318, 294.00397, 288.3746, 282.98294, 277.67044, 272.11993, 266.56924, 261.17703, 255.78465, 250.31285, 244.9995, 239.76532, 234.531, 229.5345, 224.29993, 218.9859, 213.83038, 208.59541, 203.3603, 198.04575, 192.73105, 187.41621, 182.25989, 177.02411, 171.78821, 166.47282, 161.23665, 156.07967, 150.92256, 145.5273, 140.21124, 134.4983, 129.18196, 123.865486, 118.707565, 113.62888, 108.629425, 103.78857, 99.106316, 94.18587, 89.820854, 85.13828, 80.53497, 75.534706, 70.45495, 65.93069, 61.24757, 56.40559, 51.722256, 47.35634, 42.672794, 37.989147, 33.384777, 29.018469, 24.572678, 20.285574, 15.998379, 11.711095, 6.70915, 2.9774606, NaN, NaN, 405.76584, 403.54706, 400.85275, 397.68295, 393.08664, 388.64874, 384.28998, 379.93112, 375.0174, 369.94507, 364.71408, 359.4037, 353.93463, 348.38617, 342.8376, 337.20956, 331.66064, 326.1116, 320.56238, 314.69592, 308.90857, 303.20032, 297.49194, 291.94196, 286.23325, 280.76227, 275.21182, 269.66125, 264.03122, 258.40106, 252.53282, 246.82301, 241.27167, 235.64087, 230.08922, 224.77536, 219.30273, 214.06792, 208.67432, 203.35991, 197.8867, 192.33405, 186.78122, 181.46625, 176.30978, 171.07387, 165.91716, 160.7603, 155.60333, 150.52556, 145.36833, 140.21097, 135.37086, 130.37195, 125.37291, 120.4531, 115.61253, 110.533775, 105.29618, 99.97909, 94.93963, 89.781, 84.62223, 79.93955, 75.336136, 70.81199, 66.12899, 61.366512, 56.6833, 51.9206, 47.07841, 42.39487, 37.39369, 32.471767, 27.549726, 22.78635, 18.26104, 13.894418, 9.527702, 5.160894, 2.0643733, NaN, NaN, 403.42743, 400.65387, 397.40482, 393.601, 388.13287, 382.74384, 377.03766, 371.5691, 365.94186, 360.7108, 355.55884, 350.56528, 345.65088, 340.57782, 335.5839, 330.27277, 324.80295, 320.04648, 315.21063, 309.97824, 304.5872, 299.19598, 293.64606, 288.49243, 283.41794, 278.42264, 273.5065, 268.59027, 263.6739, 258.9953, 254.3166, 249.63782, 245.11751, 240.4385, 235.68007, 230.84222, 226.16289, 221.32483, 216.40732, 211.64835, 206.80994, 201.9714, 197.2121, 192.13536, 186.74121, 181.50557, 176.19046, 170.79588, 165.55983, 160.48232, 155.32535, 150.00957, 144.6143, 139.0602, 133.74399, 128.3483, 123.031815, 118.03261, 113.03328, 108.03383, 103.431046, 98.431366, 93.51092, 88.749084, 83.82841, 79.38382, 75.17725, 71.049965, 66.763855, 62.080772, 57.71509, 53.4287, 48.983456, 44.855644, 40.489597, 36.202843, 31.83661, 27.549675, 23.421429, 19.451883, 15.323476, 10.956799, 6.6297274, 2.858352, NaN, NaN, 403.74362, 401.1286, 398.03806, 394.39273, 389.16238, 384.0904, 379.09753, 373.78754, 368.55667, 363.4842, 357.936, 352.5462, 347.077, 341.36984, 335.90033, 330.4307, 325.04016, 319.57022, 313.9416, 308.3921, 302.56494, 296.93582, 291.148, 285.4393, 279.889, 274.1007, 268.47083, 262.6822, 256.9727, 251.10443, 245.3153, 239.60533, 233.9745, 228.26422, 222.55377, 216.92247, 211.29102, 205.73874, 200.10698, 194.79236, 189.35863, 184.04373, 178.80803, 173.8102, 168.89156, 163.81415, 158.7366, 153.50026, 148.26378, 143.18585, 138.10779, 133.10896, 127.63391, 122.158714, 116.92144, 111.763374, 106.36712, 101.44687, 96.44714, 91.209206, 85.97114, 80.97103, 76.5264, 72.00229, 67.63683, 63.191902, 58.98501, 54.936783, 50.49158, 45.9669, 41.362736, 37.076008, 33.027348, 28.899221, 24.532843, 20.086979, 15.641019, 11.115568, 6.590017, 2.4613564, NaN, NaN, 403.1486, 400.69202, 397.36374, 393.7184, 388.48807, 383.81232, 378.978, 373.74725, 369.07117, 364.39502, 359.9565, 355.35938, 350.84143, 346.08557, 341.3296, 336.33572, 331.1039, 325.87195, 320.63986, 315.56622, 310.33386, 305.10138, 299.7895, 294.3982, 289.00674, 283.53586, 278.06482, 272.9901, 267.99457, 263.1575, 258.55823, 254.19673, 249.99376, 245.87, 241.74615, 237.70155, 233.41893, 229.05692, 224.61548, 220.01534, 215.25645, 210.49747, 205.73837, 200.82051, 195.7439, 190.5085, 185.19365, 180.11664, 174.56352, 169.16893, 164.17085, 159.09334, 154.09503, 149.09659, 144.09804, 139.17871, 134.33861, 129.73643, 125.372215, 121.1666, 116.92123, 112.55673, 108.112785, 103.7481, 99.46269, 95.137505, 90.89159, 86.76463, 82.677284, 78.62953, 74.34359, 70.13693, 65.850815, 61.802734, 57.635506, 53.54757, 49.022964, 44.617332, 40.29099, 35.964554, 31.717413, 27.628962, 23.738903, 19.769379, 15.6012945, 11.591915, 7.582457, 3.969908, 1.7864681, NaN, NaN, 398.94824, 396.01617, 392.37082, 388.32916, 382.5439, 376.83777, 370.97293, 365.425, 360.11465, 354.7249, 349.2558, 343.7865, 338.31708, 332.9268, 327.29852, 321.7494, 316.2794, 311.12634, 306.1317, 301.21628, 295.98358, 290.75073, 285.67636, 280.60184, 275.84436, 271.08676, 266.2498, 261.49197, 256.73407, 251.89674, 247.45581, 243.01479, 238.49437, 234.21178, 229.92908, 225.6463, 221.36343, 217.1598, 213.1147, 208.91089, 204.86565, 200.74098, 196.69557, 192.80872, 188.9218, 185.11412, 181.1874, 177.22092, 173.13538, 168.97041, 164.68637, 160.24356, 155.60231, 151.00061, 146.20047, 141.51923, 136.75853, 132.35478, 127.75258, 123.031235, 118.23043, 113.62791, 109.26334, 105.136765, 100.93075, 96.96272, 93.07398, 89.105804, 85.13755, 81.16922, 77.042076, 72.676735, 68.07319, 63.310787, 58.310143, 53.547516, 49.022915, 44.33945, 39.576496, 34.972202, 30.526579, 26.120552, 21.873213, 17.66548, 13.656146, 9.329152, 5.3196535, 2.1834567, NaN, NaN, 380.04718, 377.3526, 372.20108, 365.7021, 359.6784, 353.4168, 347.155, 340.81372, 334.71008, 328.84406, 323.29495, 317.90427, 312.3549, 306.9639, 301.4935, 295.78513, 289.918, 283.9714, 277.7075, 271.76056, 265.81345, 260.10403, 254.4738, 248.9227, 243.68867, 238.45451, 233.37883, 228.38234, 223.54436, 218.78557, 214.18529, 209.74356, 205.30173, 200.70116, 195.94183, 191.34105, 186.18489, 180.7906, 174.92018, 169.0496, 163.05986, 157.03026, 151.07983, 144.97054, 139.01976, 133.0688, 127.276375, 121.801186, 116.167145, 110.92973, 105.61282, 100.13706, 94.661156, 89.10573, 83.94699, 78.62939, 73.31164, 68.23187, 63.231358, 57.913216, 52.356796, 47.276512, 42.037334, 36.639256, 31.479195, 26.239614, 20.761728, 15.601265, 10.520068, 5.438744, 2.1040568, NaN, NaN, 299.43195, 294.43707, 288.25275, 280.48245, 273.26694, 265.49606, 257.7249, 249.79485, 241.9438, 234.17175, 226.3201, 218.54747, 210.6159, 202.92198, 195.22778, 187.69196, 180.3145, 172.77812, 165.16212, 157.62518, 150.40533, 143.26456, 136.28224, 129.37903, 122.79299, 116.12739, 109.38221, 102.79553, 96.526085, 90.09772, 83.74852, 77.79596, 72.081345, 66.36657, 60.175385, 53.58712, 47.078026, 41.124405, 34.932457, 28.502155, 21.873178, 15.045505, 8.058812, 2.9774303, NaN, NaN, 242.30055, 237.6215, 231.83203, 224.05962, 216.52484, 208.83115, 201.21649, 193.44292, 185.35173, 177.10156, 168.85107, 160.36223, 151.63503, 142.11401, 132.98929, 124.89572, 116.64313, 108.15213, 99.34334, 90.37544, 81.84367, 73.82746, 65.81093, 57.635326, 50.015057, 42.55327, 34.853054, 27.07316, 19.372362, 11.909456, 4.12869, NaN, NaN, 211.92444, 207.48267, 201.5337, 192.72893, 183.7651, 174.56291, 165.28098, 156.39531, 147.82661, 139.01953, 130.29143, 122.03905, 113.54828, 105.69202, 97.676735, 89.42304, 81.32776, 73.31152, 65.374344, 57.357487, 49.89597, 42.51356, 35.36904, 28.065498, 21.158648, 14.330955, 7.02666, 2.4216444, NaN, NaN, 196.89331, 192.21324, 186.26384, 177.22041, 168.09727, 159.13239, 150.40514, 141.99489, 133.4256, 124.7766, 115.73047, 106.84266, 98.113174, 89.46269, 81.12931, 73.11307, 65.01714, 56.762142, 48.26867, 40.171757, 32.153915, 24.135757, 16.27607, 8.25729, 2.6201377, NaN, NaN, 194.75153, 190.46803, 184.63757, 176.07007, 166.6692, 157.3869, 148.46123, 139.53517, 130.72774, 122.038956, 113.3498, 103.707985, 94.06571, 84.06584, 74.06548, 64.18369, 54.30143, 45.01405, 36.559784, 28.224253, 20.40442, 12.941561, 4.446273, NaN, NaN, 193.75993, 189.07979, 183.05098, 174.00742, 164.96347, 155.83978, 146.87436, 138.22594, 130.05324, 122.67373, 115.45266, 108.390045, 101.00975, 93.23238, 84.422966, 74.740105, 65.6124, 57.119297, 48.863987, 41.640312, 34.49577, 26.398321, 18.538727, 10.996407, 3.9301915, NaN, NaN, 185.23242, 180.59175, 174.64201, 165.83609, 156.43477, 147.033, 137.5118, 128.10916, 118.587074, 108.11227, 97.39884, 87.39914, 77.518, 67.99356, 58.825867, 50.25311, 42.27536, 34.416374, 26.795254, 19.173851, 11.194889, 3.5729034, NaN, NaN, 182.5749, 177.89452, 171.54805, 161.78996, 152.42812, 143.14519, 134.09988, 125.29223, 116.16678, 107.040924, 97.755936, 88.787994, 80.057755, 71.485886, 63.7074, 56.563633, 50.372166, 43.62484, 36.559753, 29.335653, 22.46855, 15.005772, 7.225138, 2.4613395, NaN, NaN, 176.10954, 171.82565, 165.87567, 157.46608, 149.05612, 140.56648, 131.99716, 123.66551, 115.25418, 106.60443, 97.954315, 89.70065, 82.16096, 75.097206, 67.71572, 60.492718, 53.42822, 46.680996, 40.251083, 33.900352, 27.549427, 21.357082, 15.323338, 8.813045, 3.1759155, NaN, NaN, 168.05731, 163.45593, 157.5057, 148.93707, 140.36809, 131.95744, 123.62581, 115.45254, 107.120224, 99.10501, 91.645035, 84.34351, 77.43857, 70.61277, 64.18361, 58.07175, 51.086548, 43.86296, 36.877274, 30.208893, 23.81816, 17.46692, 10.559726, 3.7316947, NaN, NaN, 160.20311, 155.44287, 149.65111, 141.79625, 134.17912, 126.085625, 117.991806, 110.135735, 102.35872, 94.740135, 87.20064, 79.89896, 72.200165, 64.26296, 56.563587, 49.340195, 42.275314, 35.52773, 28.859306, 22.031887, 14.926367, 7.4633193, 2.69953, NaN, NaN, 153.34036, 148.2626, 141.99457, 133.34596, 124.22087, 115.09538, 106.128204, 96.76383, 87.63712, 78.51, 69.064995, 59.540173, 50.173664, 40.330437, 30.883665, 21.754017, 14.5294, 6.589965, 1.8261561, NaN, NaN, 149.61137, 145.16826, 138.82079, 129.93399, 121.046814, 112.159256, 103.03323, 94.14489, 85.97044, 78.11315, 71.366745, 65.175735, 58.90516, 53.269413, 47.871655, 41.91808, 35.0911, 27.787563, 20.404379, 13.417895, 5.9150977, 1.5482635, NaN, NaN, 140.0506, 134.33774, 127.31546, 117.674324, 108.38983, 98.390686, 88.272, 78.62902, 68.985596, 59.103584, 48.74482, 39.099983, 29.573772, 20.404375, 11.472749, 3.612596, NaN, NaN, 135.76593, 130.92578, 124.41917, 115.92852, 107.59624, 98.62874, 89.89893, 80.93066, 72.27947, 64.104164, 55.452263, 46.64124, 37.353535, 28.779894, 20.285284, 11.15517, 3.2950068, NaN, NaN, 130.01324, 124.93491, 118.824875, 110.25465, 101.44598, 93.192474, 85.573555, 78.27183, 70.96984, 63.508842, 55.333183, 46.99844, 38.10767, 29.692837, 21.912777, 13.973637, 5.3990183, NaN, NaN, 133.14745, 129.25941, 122.91145, 113.944626, 105.136116, 96.48596, 88.470345, 81.32745, 74.343056, 66.961555, 59.182915, 51.007088, 43.069077, 35.051373, 27.112741, 19.65015, 11.949103, 4.0889745, NaN, NaN, 130.92569, 126.87893, 120.92765, 111.64332, 102.91408, 94.89872, 87.51796, 80.692505, 74.025566, 68.15213, 62.199146, 56.245995, 50.292667, 44.577312, 38.94118, 33.463665, 27.3509, 20.602833, 14.013328, 6.073883, 1.8261538, NaN, NaN, 124.26036, 119.4993, 112.83362, 103.66796, 93.66859, 84.14493, 74.38271, 64.262856, 53.785297, 44.021637, 34.13843, 24.96925, 16.395098, 7.5824, 1.6276592, NaN, NaN, 123.58585, 118.70575, 112.04005, 103.11243, 93.35112, 83.11315, 72.63656, 61.92131, 52.396175, 42.989666, 34.297195, 26.199764, 18.340187, 11.075764, 3.5728927, NaN, NaN, 121.80043, 116.80125, 110.01646, 100.612595, 90.49403, 80.01783, 70.49354, 61.445045, 53.229626, 45.37109, 37.15502, 28.581387, 20.483732, 12.504848, 4.4065576, NaN, NaN, 117.19798, 112.43676, 106.247, 98.62858, 91.00987, 82.67659, 73.271484, 63.984997, 54.45996, 43.98191, 34.33687, 25.167702, 16.712652, 8.376346, 2.3025367, NaN, NaN, 118.94371, 114.30155, 107.99282, 99.184074, 90.017815, 80.25589, 70.01727, 61.325954, 52.991467, 44.77571, 36.91685, 29.295855, 21.912743, 14.529363, 6.907531, 1.7864527, NaN, NaN, 120.768745, 115.76955, 109.42118, 101.08865, 92.43834, 83.62893, 75.05724, 66.96143, 58.865307, 50.05445, 41.79889, 34.495613, 27.747793, 21.396698, 15.045407, 7.741179, 2.1040418, NaN, NaN, 121.36383, 116.52335, 110.333725, 102.00124, 93.43033, 84.462234, 75.65248, 66.6836, 57.555584, 48.50654, 39.536472, 30.327856, 21.436384, 12.62392, 4.6844387, NaN, NaN, 115.80914, 111.0479, 104.69939, 96.922195, 89.70026, 81.84313, 74.303185, 66.52484, 58.587452, 50.17348, 41.44164, 32.78881, 24.215004, 16.275974, 8.257241, 2.3025336, NaN, NaN, 115.65041, 110.96851, 104.93743, 95.96984, 86.44631, 76.92233, 67.55666, 57.95243, 47.950855, 38.583855, 29.692749, 21.515764, 13.338452, 3.9698682, NaN, NaN, 109.77815, 104.77869, 98.033195, 88.66849, 78.98588, 69.46156, 59.77805, 50.332214, 41.282856, 32.391865, 24.056215, 16.196575, 7.1457057, 1.6673536, NaN, NaN, 110.73038, 106.04837, 99.85843, 91.68426, 83.033554, 74.779335, 66.52478, 58.11115, 49.776546, 42.15604, 35.090946, 28.501928, 22.150867, 15.323257, 7.939655, 2.3819287, NaN, NaN, 111.08744, 106.08801, 99.77904, 91.32709, 82.3986, 72.9935, 63.468906, 53.467606, 44.537464, 36.202312, 27.866821, 19.650076, 10.956638, 3.3346913, NaN, NaN, 107.198975, 102.43753, 96.24748, 87.596985, 79.18422, 69.9774, 60.849545, 51.80066, 42.830757, 34.257385, 25.524876, 17.347734, 9.249662, 2.818611, NaN, NaN, 103.54851, 99.104416, 92.914276, 84.18427, 74.977684, 66.405655, 57.992027, 50.05432, 42.19569, 34.89245, 27.588947, 19.808844, 11.472691, 3.4537842, NaN, NaN, 105.88951, 101.04868, 95.01733, 87.31915, 80.096886, 72.63626, 65.095985, 57.39669, 50.093994, 42.235367, 34.297054, 26.279043, 17.308027, 8.0984335, 2.6995134, NaN, NaN, 100.572495, 95.731544, 89.382576, 80.811165, 72.55687, 64.61973, 57.317295, 50.649628, 43.90236, 36.281647, 27.866785, 18.737059, 9.606927, 2.6201158, NaN, NaN, 96.9616, 92.6761, 87.04132, 79.66032, 73.07275, 66.16748, 59.420723, 52.91188, 46.40283, 39.25851, 31.955172, 24.969126, 18.141623, 10.440561, 3.3743842, NaN, NaN, 97.75518, 93.310974, 87.35876, 79.6603, 72.27903, 64.50063, 56.721947, 48.7842, 40.84615, 32.669632, 24.254623, 15.521703, 6.7090135, 1.5482534, NaN, NaN, 93.11255, 88.66824, 82.47779, 73.985466, 65.49278, 56.682247, 47.87133, 39.298183, 31.28038, 24.056149, 17.069836, 9.924497, 5.7959642, 4.7638183, NaN, NaN, 95.73146, 90.49358, 83.747635, 75.6522, 67.55645, 59.30163, 51.363983, 43.82294, 36.916687, 30.327744, 23.73859, 17.228615, 10.083283, 3.7316666, NaN, NaN, 89.1444, 84.700005, 78.74754, 70.81065, 63.270325, 55.412212, 47.315662, 39.377556, 31.597914, 23.976753, 16.4347, 8.812974, 4.605025, 2.8583035, 2.6995099, NaN, NaN, 89.144394, 84.06508, 77.47765, 68.35015, 59.301613, 50.332058, 41.838398, 33.344387, 24.453083, 15.561391, 5.9547534, 0.79397714, NaN, NaN, 87.080925, 82.47776, 76.36649, 68.50889, 61.047848, 53.0309, 44.616734, 36.281605, 28.42246, 20.563013, 13.020835, 6.9868927, 4.446232, 3.8904583, NaN, NaN, 90.89036, 85.573, 78.98562, 70.0963, 60.968468, 51.602097, 42.314682, 33.423767, 24.532467, 15.6407795, 6.5899158, 1.587951, NaN, NaN, 89.937996, 85.89044, 80.255486, 73.58857, 67.23893, 60.333466, 53.427773, 46.442467, 39.695072, 32.86807, 25.88206, 18.34008, 11.19479, 6.5105195, 4.922607, NaN, NaN, 83.94599, 78.866554, 72.437706, 63.230606, 54.023094, 45.21207, 36.2419, 27.82705, 19.570631, 11.075698, 2.8186038, NaN, NaN, 87.47771, 82.71582, 76.5252, 68.112, 59.777832, 51.60208, 43.267242, 35.09083, 27.072868, 19.05459, 10.8772135, 5.478377, 3.572871, 3.414078, NaN, NaN, 83.78725, 79.50147, 73.628235, 64.73868, 55.68999, 46.482143, 37.591415, 28.779686, 19.808796, 10.599335, 2.6598096, NaN, NaN, 83.11265, 78.43002, 72.31864, 64.22276, 56.60282, 48.823837, 41.04456, 33.423756, 24.9294, 15.878949, 7.9396286, 4.049249, 2.2231271, NaN, NaN, 87.47772, 82.7952, 76.84268, 68.66761, 60.650963, 52.87213, 45.489906, 39.06001, 33.26499, 25.802671, 17.069824, 8.6541815, 2.937699, NaN, NaN, 92.239525, 87.39838, 81.128525, 72.79488, 64.30216, 55.809082, 47.712547, 40.4889, 33.18561, 25.008797, 16.67287, 8.654183, 3.9698544, 2.2231278, NaN, NaN, 91.84273, 87.1603, 81.12854, 73.11238, 65.0959, 56.84098, 48.34759, 39.377556, 30.88344, 22.706532, 14.76747, 6.4311266, 1.508554, NaN, NaN, 98.07259, 92.59669, 85.21589, 75.92999, 67.51676, 60.21444, 52.59434, 44.8152, 37.829597, 33.622242, 27.668293, 18.538567, 10.12298, 3.771365, 1.7864447, NaN, NaN, 92.953835, 87.71589, 81.525406, 72.080605, 63.032227, 54.30096, 45.56932, 36.281624, 26.91412, 18.101921, 9.765709, 2.8583045, NaN, NaN, 102.11995, 97.040955, 90.45394, 82.120674, 74.10454, 65.77061, 57.11883, 48.784206, 40.846153, 32.74902, 25.048512, 17.506493, 9.09086, 2.8980036, NaN, NaN, 103.905525, 99.46145, 93.430046, 85.33499, 77.63646, 69.85826, 62.476643, 55.729763, 49.53832, 43.10854, 35.170265, 26.755356, 18.657665, 12.0681305, 4.446236, NaN, NaN, 103.98491, 99.54083, 93.985596, 86.20802, 78.350784, 69.30268, 59.857304, 51.046516, 43.505455, 37.234253, 30.7247, 23.738611, 15.6407995, 7.383877, 2.3819249, NaN, NaN, 101.28676, 96.287094, 90.17624, 82.160416, 74.30302, 65.651596, 57.317314, 49.06207, 40.80649, 32.94751, 25.961493, 18.657675, 10.480265, 2.8583074, NaN, NaN, 108.349594, 103.42946, 97.08073, 89.2239, 81.84297, 74.22367, 66.60408, 58.031708, 49.06208, 40.64774, 31.994892, 23.42107, 14.60871, 5.3989925, NaN, NaN, 111.96029, 107.27831, 100.9297, 92.04131, 83.152534, 75.37454, 68.231224, 60.770164, 52.435677, 44.02147, 35.6863, 27.112629, 19.094334, 11.552087, 3.8507679, NaN, NaN, 113.983864, 109.301926, 103.03274, 94.303154, 85.97003, 77.080986, 67.7947, 58.58737, 49.697144, 41.044674, 32.23307, 23.73864, 15.482034, 7.939651, 2.2231333, NaN, NaN, 121.1653, 116.72159, 110.849396, 103.31052, 96.247536, 89.02557, 81.4859, 74.18405, 66.723206, 58.547703, 49.73685, 40.76685, 32.51093, 25.207336, 18.53861, 11.313912, 4.485942, NaN, NaN, 117.316765, 112.71426, 106.683235, 99.382286, 92.31916, 84.62087, 77.23977, 70.09651, 62.39739, 54.38047, 44.855007, 35.3291, 27.07296, 19.927952, 13.100266, 5.9547706, 1.4291607, NaN, NaN, 122.990425, 118.11031, 111.801704, 102.8741, 93.946106, 85.01772, 76.32705, 68.2313, 59.89711, 50.371902, 39.298294, 30.367525, 24.175297, 17.387447, 8.932093, 2.620121, NaN, NaN, 124.617134, 119.73706, 113.4285, 105.33421, 97.23961, 88.90659, 79.97799, 70.81088, 62.59585, 54.618626, 45.688522, 37.710636, 31.280474, 22.349354, 11.631495, 3.294996, NaN, NaN, 124.73618, 119.61806, 113.071434, 104.38195, 95.6921, 85.69236, 74.858765, 64.381775, 55.452095, 47.712727, 41.282875, 33.185734, 23.897448, 14.966004, 6.272358, 1.9849441, NaN, NaN, 126.680275, 122.07798, 116.12658, 107.397545, 98.27134, 89.22409, 80.81138, 72.95391, 65.01677, 56.92057, 49.220943, 41.362267, 33.26513, 25.405836, 18.181374, 10.87726, 3.8110766, NaN, NaN, 127.83087, 123.06989, 116.88046, 108.23081, 99.104645, 89.81934, 80.374886, 71.48558, 63.31026, 55.45212, 47.27616, 38.464806, 29.732462, 22.428759, 15.442365, 7.423596, 2.3422332, NaN, NaN, 128.78308, 124.02213, 118.070786, 109.73861, 101.247375, 92.91451, 84.74004, 76.40652, 67.75516, 59.10343, 50.927616, 43.30714, 35.924538, 28.382893, 20.602798, 12.266656, 4.5653462, NaN, NaN, 134.93253, 130.40976, 124.458595, 115.17443, 105.73114, 97.3191, 89.30353, 81.60512, 73.35082, 64.85808, 56.60311, 48.98285, 41.67983, 34.37655, 27.390558, 20.086767, 11.988782, 4.843235, 0.7939808, NaN, NaN, 136.4798, 131.56033, 125.05375, 115.531555, 106.64377, 97.596886, 89.18451, 80.77178, 72.6762, 64.73904, 56.72219, 49.02255, 41.71953, 34.654404, 27.112707, 20.36464, 13.219382, 5.6768966, 1.3894647, NaN, NaN, 139.05855, 134.77391, 128.58482, 120.37209, 112.159035, 103.58854, 94.06534, 84.7798, 75.851, 67.39804, 59.182858, 50.61014, 42.751507, 37.15502, 30.724827, 20.7219, 10.956669, 3.5728912, NaN, NaN, 142.82741, 138.38416, 132.27454, 123.86357, 115.29356, 106.80254, 98.31118, 89.89883, 81.3274, 72.67624, 64.58033, 57.277855, 50.133884, 41.9577, 33.939957, 26.715784, 19.729527, 12.98121, 6.3120675, 2.262839, NaN, NaN, 152.50708, 148.3814, 142.90681, 135.92451, 129.18002, 121.56245, 113.78587, 106.4058, 98.78738, 90.85122, 82.91476, 75.13673, 67.19965, 59.897274, 53.547165, 46.6412, 39.496857, 32.907963, 26.398241, 19.729534, 12.901822, 6.232674, 2.104045, NaN, NaN, 156.31538, 151.47572, 145.2078, 137.35277, 129.81485, 121.64183, 113.389145, 105.05676, 97.2002, 89.81953, 82.51795, 74.89864, 66.644066, 58.309784, 50.05454, 42.75155, 35.686447, 27.986006, 20.126493, 12.743039, 5.2402244, 1.3894665, NaN, NaN, 164.48706, 159.96494, 153.7766, 145.52519, 137.5115, 129.49748, 121.562515, 113.23046, 104.659996, 96.16854, 87.83546, 79.66077, 71.961975, 64.58039, 57.277912, 50.133934, 42.83094, 36.4803, 30.447012, 23.77843, 16.75237, 9.448189, 3.6522927, NaN, NaN, 171.54778, 166.78781, 160.52034, 152.42789, 144.96985, 137.03548, 128.9421, 120.61034, 112.51631, 104.739395, 97.1209, 89.42277, 81.48624, 73.5494, 66.0885, 58.944824, 52.118416, 44.97425, 37.512306, 30.129475, 22.547903, 15.640887, 9.130612, 3.1759114, NaN, NaN, 178.05296, 173.29314, 167.10521, 159.01302, 151.39653, 143.62108, 135.92468, 127.83126, 119.658165, 111.40538, 103.072914, 94.97819, 87.35933, 79.81956, 71.96203, 64.02482, 56.484188, 49.498936, 42.513443, 35.13079, 27.350933, 20.523466, 14.17213, 7.1060367, 2.1040478, NaN, NaN, 186.18414, 181.42451, 174.84016, 166.27226, 157.30733, 148.50067, 139.77298, 131.04492, 122.15778, 113.42898, 104.77915, 96.20833, 87.87524, 79.46244, 70.73181, 61.84206, 53.50757, 44.934597, 37.075726, 30.248579, 23.421207, 15.958469, 9.051225, 3.4141057, NaN, NaN, 191.81631, 186.7395, 180.15532, 171.19098, 161.35356, 152.7851, 144.05759, 134.77428, 126.363396, 118.269585, 110.49288, 102.874596, 94.93858, 87.08162, 79.06563, 71.20806, 62.953323, 55.015762, 47.236652, 40.09231, 33.424038, 26.43799, 18.816578, 11.988821, 5.002044, 1.0321778, NaN, NaN, 203.47675, 199.03479, 193.00627, 185.5497, 178.4895, 171.0324, 163.33702, 155.80003, 147.78673, 139.69376, 131.52112, 123.427505, 115.49229, 107.556755, 99.70027, 91.76413, 83.82768, 76.129036, 68.35072, 60.730865, 53.428238, 46.20473, 39.2985, 32.94774, 25.882284, 18.816587, 12.782764, 6.1929917, 2.1437492, NaN, NaN, 231.43518, 226.67659, 220.173, 211.44835, 203.27856, 195.26709, 187.33464, 179.48122, 171.86548, 164.17014, 156.0778, 147.74713, 139.09875, 130.84674, 123.070496, 115.690735, 107.91392, 100.05745, 92.359406, 84.42297, 76.68466, 68.906364, 61.0484, 53.34889, 45.56971, 38.584072, 31.995125, 25.802912, 19.451727, 13.735493, 8.257285, 3.1759186, NaN, NaN, 308.7868, 303.9507, 297.60812, 289.1246, 280.79932, 272.4737, 264.14774, 255.58354, 247.2569, 238.77132, 230.20605, 221.71976, 213.15381, 204.66681, 196.25877, 187.69176, 179.12437, 170.87396, 162.62321, 154.21347, 145.92238, 137.74998, 129.89465, 122.27708, 114.65922, 106.961716, 99.1052, 90.85158, 82.75635, 75.05765, 67.5174, 60.29438, 53.071106, 46.1651, 39.417625, 32.749317, 26.398344, 19.809, 13.7752, 7.106055, 2.4216442, NaN, NaN, 382.66214, 378.06555, 372.12152, 363.48254, 354.76395, 345.88644, 337.1671, 328.7645, 320.4408, 312.19608, 304.34738, 296.4984, 288.56985, 280.7996, 273.1083, 265.02023, 256.9319, 248.76389, 240.59557, 232.26831, 223.70279, 214.74033, 205.85678, 197.29015, 188.80249, 180.79045, 173.01608, 165.79677, 158.73589, 151.99211, 145.01009, 137.47241, 129.77576, 121.92011, 114.381584, 107.318924, 100.73218, 93.986496, 87.002495, 79.78015, 72.31945, 64.7791, 57.63535, 50.491352, 43.267723, 36.52015, 30.010511, 23.659449, 17.546362, 11.830066, 6.034213, 2.064356, NaN, NaN, 488.75232, 484.4749, 479.00922, 471.08768, 463.4827, 455.719, 448.43036, 441.2207, 434.01077, 426.87985, 419.51096, 412.3003, 405.0101, 397.4027, 389.55728, 381.7908, 373.8655, 365.9399, 358.01404, 349.85004, 341.68573, 333.83817, 326.46594, 318.93494, 311.40363, 303.87204, 296.1816, 288.57016, 281.03775, 273.66364, 266.36856, 259.15253, 251.69832, 244.48177, 237.10635, 229.65135, 221.95815, 214.34396, 206.80882, 199.11476, 191.61873, 184.24141, 177.18115, 170.27931, 163.61523, 156.55426, 149.81041, 142.90765, 136.084, 129.57751, 123.22954, 117.04006, 110.77104, 104.58119, 98.39116, 91.88348, 85.058136, 78.3913, 71.96236, 66.00945, 59.977, 54.02375, 47.752804, 41.64043, 35.44849, 29.891462, 24.096115, 18.459387, 12.663716, 6.8678803, 2.501047, NaN, NaN, 500.436, 495.9212, 489.98056, 481.66336, 473.02896, 464.63187, 456.15518, 447.91586, 439.7554, 431.6739, 423.43356, 415.66837, 407.74435, 399.97858, 391.97473, 383.73282, 375.56985, 367.4858, 359.40146, 351.31677, 343.1525, 335.14645, 327.45718, 320.00546, 312.3949, 304.46695, 296.61795, 288.45154, 280.36407, 272.3556, 264.58466, 256.81345, 249.12126, 241.34947, 233.8153, 226.28088, 218.74617, 211.13187, 203.75523, 196.37834, 189.15984, 181.94109, 174.8014, 167.58214, 160.5213, 153.69823, 146.7956, 139.57533, 132.19614, 124.57862, 116.80212, 109.025314, 101.4863, 94.34382, 87.51855, 80.45495, 73.15299, 66.16827, 59.659557, 53.46816, 47.67347, 41.958004, 36.401146, 31.161686, 25.92209, 20.44419, 14.807354, 8.9321785, 3.453822, NaN, NaN, 498.53568, 493.94165, 488.00095, 480.39658, 473.02957, 465.2662, 457.34412, 449.3425, 441.4198, 433.41754, 425.57346, 417.49136, 409.64667, 401.8017, 394.1149, 386.6656, 379.21597, 371.7661, 364.23672, 356.94482, 349.53378, 342.08286, 334.4731, 326.94235, 319.1735, 311.24576, 303.47632, 295.548, 287.93652, 280.48337, 273.1885, 266.052, 258.9945, 251.7782, 244.32372, 236.78966, 229.17603, 221.24484, 213.63062, 206.17474, 198.79794, 191.57951, 184.44016, 177.14189, 169.76402, 162.22723, 154.53148, 146.9148, 139.53584, 132.15663, 125.253265, 118.429016, 111.52518, 104.462395, 97.161285, 90.3361, 83.986885, 77.558105, 71.36723, 65.4143, 59.659634, 54.262005, 48.943615, 43.30756, 37.830116, 32.74946, 27.906837, 23.540443, 19.015171, 14.0928335, 8.614608, 3.4538264, NaN, NaN, 499.68497, 495.48697, 489.94235, 482.65488, 475.5256, 468.3961, 460.94943, 453.66095, 446.13452, 438.60782, 430.9224, 423.4744, 415.94687, 408.41907, 400.7325, 393.0457, 385.4378, 377.82965, 370.30045, 363.00876, 355.75647, 348.46426, 341.01328, 333.562, 326.11047, 318.42087, 311.04807, 303.5957, 296.1431, 288.92807, 281.55423, 274.2594, 266.80573, 259.51038, 251.89755, 244.12584, 236.11592, 228.34361, 220.33307, 212.08427, 204.31107, 196.77553, 189.557, 182.25891, 174.96056, 167.50328, 160.04573, 152.42923, 144.49507, 136.95734, 129.97476, 123.15066, 116.326324, 109.10499, 101.80403, 94.344086, 87.67753, 81.32822, 74.81998, 68.31152, 61.92193, 56.60373, 51.206013, 45.252483, 39.06063, 33.344906, 28.343515, 23.977123, 18.896114, 13.65619, 7.2251906, 2.7789497, NaN, NaN, 500.04214, 495.52734, 489.66586, 482.06155, 475.09067, 467.80267, 460.59363, 453.22592, 445.7787, 438.3312, 430.96268, 423.43542, 416.06638, 408.53857, 401.169, 393.5614, 385.87427, 378.34537, 371.1332, 364.00006, 356.94595, 349.8123, 342.6784, 335.2272, 327.85498, 320.32397, 312.63412, 305.10254, 297.4914, 289.95926, 282.34756, 274.81488, 267.4405, 260.06586, 252.69095, 245.15718, 237.70244, 230.0888, 222.47488, 214.86069, 207.12723, 199.59178, 192.45268, 185.39265, 178.17374, 170.95456, 163.73512, 156.4361, 149.21616, 141.99597, 134.9342, 127.87221, 120.80997, 114.14426, 107.7164, 100.89155, 94.14583, 87.24115, 80.733086, 74.304184, 67.875084, 61.366398, 55.095646, 49.14222, 43.18862, 37.155464, 30.963354, 24.850449, 19.13432, 13.894393, 7.9397683, 3.0171483, NaN, NaN, 498.26065, 493.6666, 487.72586, 479.4085, 471.4077, 463.64426, 455.72205, 447.72034, 439.63907, 431.5575, 423.31714, 414.8387, 406.35995, 398.19785, 389.71838, 381.31784, 372.59995, 364.1987, 355.95563, 347.71225, 339.58743, 331.34338, 323.4161, 315.72635, 308.1949, 300.4253, 292.73468, 285.36093, 277.59045, 269.9783, 262.44516, 254.99101, 247.53662, 240.16125, 232.62701, 225.1718, 217.24043, 209.62604, 202.09067, 194.47571, 186.78113, 178.84827, 171.07378, 163.37833, 155.84126, 148.62129, 141.32172, 134.0219, 126.5631, 119.73886, 113.23182, 106.56586, 99.89967, 93.23328, 86.64603, 80.45541, 74.50271, 68.62921, 63.073048, 57.119846, 51.285538, 45.728905, 40.48965, 35.32965, 30.090134, 25.644377, 21.516087, 17.387714, 13.179864, 8.495552, 3.5729387, NaN, NaN, 499.9643, 495.5287, 489.7464, 481.90442, 474.379, 466.77408, 459.08966, 451.40497, 443.7992, 435.95547, 428.11142, 420.0294, 412.10553, 404.02286, 395.93985, 387.93582, 380.1692, 372.2438, 364.31808, 356.23355, 348.18832, 340.34094, 332.65182, 324.88312, 317.19342, 309.50342, 302.051, 294.36044, 286.19385, 278.50272, 270.89056, 263.11954, 255.11032, 247.2594, 239.48747, 231.79459, 223.86345, 215.8527, 207.92096, 199.98892, 191.97723, 184.04457, 176.27026, 168.89233, 161.67282, 154.53238, 147.55038, 140.25076, 132.79219, 125.65074, 118.90582, 111.92261, 104.54236, 97.16185, 90.257256, 83.74927, 77.24107, 70.49456, 64.22407, 58.112137, 52.238163, 46.52278, 40.80724, 34.456455, 28.502413, 22.86576, 18.022879, 13.021093, 7.0664277, 2.5407662, NaN, NaN, 498.65808, 493.9848, 487.96484, 479.48907, 471.17136, 463.01178, 454.9311, 446.92932, 438.92725, 430.92484, 422.92212, 414.99835, 407.39124, 399.8631, 392.57242, 385.2815, 378.06955, 370.69882, 363.2486, 355.71884, 348.34735, 340.81705, 333.28644, 325.67633, 317.90735, 310.37595, 302.68567, 294.99515, 287.3043, 279.77176, 272.23895, 264.70587, 257.4104, 249.95605, 242.34285, 235.04659, 227.75008, 220.61192, 213.23557, 206.09692, 198.99768, 191.54123, 184.3225, 177.1035, 169.9636, 162.90277, 155.8417, 148.7804, 141.87753, 135.21248, 128.62656, 122.11978, 115.53344, 108.946884, 102.67756, 96.56677, 90.69389, 84.90021, 78.947624, 72.75675, 66.52601, 60.41414, 54.460842, 48.427994, 42.95065, 37.87008, 33.18632, 28.740618, 24.85055, 20.722233, 15.958687, 10.639263, 4.605122, 1.1909897, NaN, NaN, 498.5795, 493.90622, 488.12387, 480.44025, 473.07318, 465.62665, 458.33826, 451.04965, 443.91922, 436.3924, 429.02377, 421.81335, 414.68192, 407.39175, 400.33908, 393.28613, 386.47073, 379.57584, 372.75995, 365.7061, 358.65198, 351.67688, 344.93936, 337.88452, 331.06726, 324.09125, 317.115, 310.21777, 303.3203, 296.6605, 289.92117, 283.3402, 276.759, 270.25693, 263.67532, 257.17282, 250.43219, 244.00858, 237.58475, 230.92279, 224.3796, 217.79652, 211.05461, 204.23315, 197.49078, 190.51024, 183.29144, 176.15175, 168.85312, 161.63358, 154.49312, 147.19373, 140.13211, 133.54634, 127.35712, 121.08835, 114.58132, 108.15345, 101.963455, 96.01135, 90.21782, 84.66222, 79.02709, 73.31245, 67.756386, 62.120796, 56.485054, 50.92854, 45.451252, 40.132587, 35.051945, 29.971172, 25.287226, 20.682564, 16.554157, 12.266878, 7.5031295, 3.612652, NaN, NaN, 499.7681, 495.41168, 489.78778, 482.26263, 475.05408, 467.36993, 460.0024, 452.6346, 445.34576, 437.89822, 430.3712, 422.9231, 415.55396, 408.34308, 401.13193, 393.76202, 386.3126, 378.8629, 371.1752, 363.64572, 356.23483, 348.7841, 341.41232, 334.04028, 326.8265, 319.61252, 312.39825, 305.34232, 298.04828, 290.91254, 283.77658, 276.71964, 269.74176, 262.68436, 255.62671, 248.72742, 241.7486, 234.53162, 227.31436, 220.09688, 212.95844, 205.9784, 198.9188, 192.09694, 185.35417, 179.00783, 172.50264, 165.91791, 159.17427, 152.11307, 145.13095, 138.70404, 132.03886, 125.53218, 119.42205, 113.391106, 107.28062, 101.09059, 94.97974, 88.70997, 82.12254, 75.61427, 69.185165, 62.83524, 56.723244, 50.84921, 45.292534, 40.05324, 34.97259, 30.05059, 25.28725, 20.12684, 15.045695, 9.567444, 4.803627, 1.8658851, NaN, NaN, 499.8478, 495.41217, 489.70908, 481.5502, 473.4702, 465.7068, 457.86386, 450.17908, 441.9394, 434.09555, 426.33066, 418.56546, 410.95844, 403.11343, 395.7436, 388.215, 380.84464, 373.15698, 365.62756, 358.17712, 350.56787, 342.8791, 335.19003, 327.57996, 319.73175, 311.804, 303.71735, 296.0268, 288.1774, 279.93124, 272.16052, 264.23093, 256.0631, 247.81567, 239.72652, 231.47842, 223.23, 215.21918, 207.20807, 199.35527, 192.09712, 184.71973, 177.58006, 170.20215, 162.66528, 155.04881, 147.59074, 140.37044, 133.30856, 126.563866, 120.215706, 113.39122, 106.5665, 100.059, 93.71002, 87.67831, 81.646416, 75.69372, 69.5821, 63.629055, 58.152096, 52.516235, 46.800835, 41.64096, 36.08403, 30.685724, 25.684225, 20.761997, 15.760255, 10.678995, 5.5182123, 2.3422809, NaN, NaN, 499.53156, 494.85828, 488.67987, 480.2041, 471.88638, 463.806, 455.40842, 447.32742, 439.32532, 430.8475, 422.84476, 414.8417, 406.91757, 399.0724, 391.3854, 383.6189, 376.1691, 368.63977, 360.6346, 353.02545, 345.45566, 337.76666, 329.8396, 322.07074, 314.3016, 306.61148, 298.84174, 290.91318, 282.7464, 274.6586, 266.4119, 258.79926, 251.18636, 243.57315, 236.2769, 229.05971, 221.525, 214.22797, 206.53407, 198.8399, 191.10577, 183.72833, 176.19196, 168.97266, 161.59442, 154.05724, 146.67847, 139.06139, 131.60272, 124.3025, 117.00201, 110.17741, 103.43193, 97.003685, 90.97206, 85.17836, 79.622604, 73.98733, 68.3519, 62.875057, 57.23932, 51.682808, 46.205524, 40.569324, 35.25052, 30.249125, 25.40639, 20.325363, 15.482394, 10.63931, 6.034303, 2.461382, NaN, NaN, 501.94794, 497.51233, 491.65085, 483.33362, 475.01602, 466.6189, 458.2214, 449.82358, 441.50464, 433.18536, 424.86575, 416.38736, 407.67084, 399.1917, 390.7915, 382.15317, 373.8315, 365.66803, 357.742, 349.73642, 342.04758, 334.4377, 326.8276, 319.1379, 311.44794, 303.51984, 295.74997, 287.82126, 280.05084, 272.3594, 264.90558, 257.29288, 249.60059, 242.22523, 234.77031, 227.31511, 219.93896, 212.40392, 204.70995, 197.17435, 189.87643, 182.41962, 174.96252, 167.58449, 160.28554, 152.90698, 145.76619, 139.10123, 132.27734, 125.53259, 118.94633, 112.35985, 105.93187, 99.42434, 93.154686, 87.20231, 81.4085, 75.69389, 69.979126, 64.10545, 58.668182, 53.032322, 47.31692, 41.680748, 36.282578, 31.281204, 26.20032, 21.039915, 16.117563, 11.512674, 5.557924, 1.9849901, NaN, NaN, 499.37424, 494.78015, 488.76016, 480.68045, 473.07568, 465.31223, 457.5485, 449.62598, 441.86163, 434.17624, 426.56976, 418.6461, 410.64285, 402.6393, 394.79395, 387.10678, 379.4986, 371.65234, 363.80582, 355.8797, 348.23074, 340.1455, 332.377, 324.529, 316.8392, 309.22842, 301.3795, 293.451, 285.76004, 278.06882, 270.3773, 262.7648, 254.99341, 247.30103, 239.68767, 232.15334, 224.69803, 217.00452, 209.2314, 201.61662, 194.23955, 186.8622, 179.64325, 172.50339, 165.44261, 158.46092, 151.47899, 144.4175, 137.51443, 130.8492, 124.342445, 117.994194, 111.88382, 105.931984, 100.37678, 95.05951, 89.50401, 84.18646, 78.63067, 72.91598, 67.63768, 62.478317, 56.921936, 51.44478, 45.888096, 40.807568, 36.044456, 31.440014, 26.914854, 22.15142, 17.387877, 12.227245, 6.6694975, 2.5407865, NaN, NaN, 500.00836, 495.65192, 490.02798, 482.58203, 475.29422, 467.84772, 460.48016, 452.9539, 445.5858, 437.9005, 430.45267, 423.00455, 415.2392, 407.47354, 399.7076, 392.02063, 384.2541, 376.40802, 368.4824, 360.87354, 353.02655, 345.25858, 337.411, 329.64243, 321.95285, 314.1837, 306.33493, 298.5652, 290.87442, 283.42126, 275.88852, 268.1969, 260.6636, 252.97144, 245.27898, 237.66554, 230.21043, 222.993, 215.77531, 208.55737, 201.25986, 193.88277, 186.58473, 179.28644, 172.14655, 164.7684, 157.46933, 150.17, 143.18779, 136.04665, 128.90524, 122.16037, 115.7327, 108.98738, 101.92441, 95.33737, 89.06758, 83.19444, 77.63862, 71.6064, 65.69308, 60.057396, 54.262806, 48.626812, 43.308197, 38.06883, 32.67055, 27.430912, 22.34992, 17.348196, 12.50514, 8.21775, 4.009668, 1.707096, NaN, NaN, 501.43463, 497.07822, 491.37512, 484.16684, 477.0375, 469.43262, 461.90665, 454.3012, 446.93317, 439.1687, 431.5624, 423.87662, 415.87357, 407.8702, 399.94577, 391.86255, 383.69977, 375.14038, 366.73914, 358.33755, 350.05453, 341.89008, 333.7253, 325.5602, 317.55334, 309.86328, 302.4108, 295.1959, 287.74286, 280.36887, 272.91528, 265.30286, 257.45227, 249.83926, 242.14667, 234.37448, 226.83994, 218.98785, 211.45274, 203.91737, 196.54036, 189.40106, 182.02353, 174.8044, 167.82301, 160.76205, 153.70085, 146.63942, 139.57773, 132.43645, 125.136215, 117.75637, 110.45562, 103.55141, 96.726326, 89.980385, 83.23422, 77.04343, 70.931816, 64.8994, 59.025562, 52.913414, 47.118614, 41.403034, 35.687294, 30.288948, 24.572897, 18.936079, 13.378502, 8.058965, 3.2950833, NaN, NaN, 502.30646, 497.87085, 492.08856, 484.00894, 475.69135, 467.53186, 459.13437, 450.49887, 442.02148, 433.62296, 425.38257, 416.98337, 408.34613, 399.94623, 391.7045, 383.30392, 375.06152, 366.58102, 358.4172, 350.33237, 342.32645, 334.32022, 326.47223, 318.3861, 310.45825, 302.53006, 294.60156, 286.59348, 278.98157, 271.21075, 263.36035, 255.66827, 248.05519, 240.44183, 232.8282, 225.05565, 217.52075, 210.06491, 202.68811, 195.23172, 187.81473, 180.35779, 172.90059, 165.44313, 158.30273, 151.32079, 144.3386, 137.19748, 130.21481, 123.31126, 116.32812, 109.10666, 102.361115, 95.2979, 88.86936, 82.44063, 75.85295, 69.82067, 64.10572, 58.390606, 52.91347, 47.59496, 42.355686, 37.19567, 31.797358, 26.795855, 21.794228, 16.792479, 11.949399, 7.026808, 2.8980913, NaN, NaN, 498.50497, 493.83163, 487.8116, 479.89023, 472.0478, 464.04657, 456.1243, 448.4394, 440.35806, 432.2764, 424.3529, 416.34985, 408.26724, 400.34283, 392.25958, 384.2553, 376.17145, 368.2458, 360.16132, 352.0765, 343.99136, 335.7474, 327.58237, 319.49628, 311.64774, 303.71957, 295.71185, 287.94168, 280.09192, 272.55902, 264.86728, 257.17523, 249.4829, 241.71097, 233.46289, 225.69037, 217.99686, 210.30305, 202.6883, 195.15257, 187.61658, 180.0803, 172.6231, 165.1656, 157.78719, 150.17047, 142.71216, 135.25359, 127.71539, 120.811745, 113.828514, 107.08312, 100.654945, 94.38531, 88.2742, 82.08355, 75.89271, 70.17792, 64.304214, 58.430347, 52.51662, 46.80118, 41.40312, 36.084297, 30.844728, 25.763805, 20.682756, 15.601583, 10.361489, 5.518253, 2.5010972, NaN, NaN, 499.0993, 494.5844, 488.5644, 480.16776, 471.77075, 463.29422, 454.89655, 446.4193, 437.7833, 429.38458, 420.9063, 412.34842, 403.9487, 395.62787, 387.38593, 379.22293, 371.21814, 363.2923, 355.28687, 347.43967, 339.59216, 331.90292, 323.97556, 315.8893, 307.88205, 299.87448, 291.8666, 284.17557, 276.32565, 268.63403, 260.86282, 253.40854, 246.1919, 238.97499, 231.91646, 224.93701, 217.9573, 210.81874, 203.75925, 196.77882, 190.11548, 183.29326, 176.55016, 169.88615, 162.98392, 156.00212, 149.02008, 141.95847, 135.0553, 127.99319, 120.93084, 113.94761, 107.20222, 100.77405, 94.34567, 87.9171, 81.647064, 75.535576, 69.82077, 64.10581, 58.192245, 52.7151, 47.555336, 41.99852, 36.7591, 31.837097, 26.914978, 21.913347, 16.911594, 11.989115, 6.7489257, 2.9377952, NaN, NaN, 498.22842, 493.4759, 487.37662, 478.9007, 470.6621, 462.5816, 454.50082, 446.7366, 439.05136, 431.3658, 423.7592, 416.23157, 408.6244, 401.01697, 393.40924, 385.8805, 378.19296, 370.66367, 363.0548, 355.52496, 347.79666, 340.1077, 332.41846, 324.57037, 316.72202, 309.0319, 301.18292, 293.25436, 285.4841, 277.79282, 270.10123, 262.33008, 254.24142, 245.91454, 237.98384, 230.05286, 222.51813, 214.90381, 207.44785, 199.99161, 192.81274, 185.59396, 178.5336, 171.71098, 164.72948, 157.74773, 151.00377, 144.41827, 137.59453, 130.61186, 123.78765, 117.20129, 110.29728, 103.71048, 97.52029, 91.17117, 85.2187, 79.42479, 73.63072, 67.677734, 61.526142, 55.414047, 49.619297, 44.062534, 38.505623, 32.948555, 27.629509, 22.310326, 16.991003, 12.465499, 7.939896, 3.5729914, NaN, NaN, 499.93198, 495.3379, 489.15945, 480.52518, 471.6529, 462.701, 453.82794, 444.9545, 436.23914, 427.44418, 418.64883, 410.40784, 402.16647, 393.76633, 385.44507, 376.80643, 368.56375, 360.2415, 351.99814, 343.75446, 335.62933, 327.54355, 319.69528, 311.76743, 303.83926, 296.14868, 288.45776, 280.92517, 273.47162, 266.09705, 258.72223, 251.26785, 244.13043, 236.99275, 229.77553, 222.55803, 215.26097, 207.96365, 200.58676, 192.89229, 185.31653, 177.70082, 169.92616, 162.30988, 154.85199, 147.39384, 140.01477, 132.87347, 125.731926, 118.98691, 112.5591, 106.369156, 99.94095, 93.433174, 86.92519, 80.25826, 73.59112, 67.24126, 60.891197, 54.85846, 49.26214, 43.70536, 38.14843, 32.829514, 27.351677, 22.032478, 16.951324, 12.1082325, 7.10623, 3.1362994, NaN, NaN, 498.74445, 493.99188, 488.13025, 480.3673, 473.00015, 465.47427, 457.86893, 449.86716, 442.18198, 434.25882, 426.1769, 418.49084, 411.04224, 403.51413, 395.98572, 388.45706, 380.84885, 373.47815, 366.0279, 358.41888, 351.16626, 343.55667, 336.0261, 328.5745, 321.12265, 313.90836, 306.53525, 299.24115, 292.0261, 284.89008, 277.7538, 270.61728, 263.48053, 256.26422, 249.04765, 242.06874, 234.85168, 227.47574, 220.25816, 213.11964, 205.90157, 198.60391, 191.38531, 184.32513, 177.2647, 170.44203, 163.69847, 157.03404, 150.29004, 143.78386, 137.27747, 130.92957, 124.58147, 118.23318, 112.122765, 105.85345, 99.42521, 92.99678, 86.726875, 80.45678, 74.424614, 68.47164, 62.677246, 57.200203, 51.64363, 45.848763, 40.37127, 35.052402, 29.733397, 24.414255, 19.094975, 14.331323, 9.885147, 4.6448874, 1.9453076, NaN, NaN, 498.9825, 494.4676, 488.52673, 480.52615, 472.92133, 464.92014, 456.83942, 448.99603, 441.2316, 433.70456, 426.09802, 418.2535, 410.25018, 402.08804, 393.68787, 385.12885, 376.88647, 368.48523, 360.00443, 351.6818, 343.43808, 335.19403, 327.02893, 318.86353, 310.77707, 302.76956, 294.60318, 286.1986, 277.873, 269.7849, 261.61722, 253.2906, 245.20157, 237.19151, 229.26047, 221.40843, 213.6354, 205.86209, 198.08847, 190.39389, 182.77837, 175.0832, 167.2291, 159.29535, 151.12326, 143.10954, 135.25421, 127.39857, 119.78069, 112.479965, 105.3377, 98.19518, 91.5286, 84.78245, 78.353546, 72.241936, 66.36827, 60.335682, 54.382294, 48.82564, 43.427605, 38.108814, 32.869274, 27.470818, 22.151611, 17.943785, 13.815266, 8.495705, 3.5730028, NaN, NaN, 500.5671, 496.21066, 490.42828, 483.1407, 476.01126, 468.40628, 460.56335, 453.11624, 445.5104, 437.9043, 430.0602, 422.13657, 414.45035, 406.68463, 398.99783, 390.99374, 382.91013, 375.22244, 367.5345, 360.00476, 352.23697, 344.70667, 337.17612, 329.48672, 321.95563, 314.26566, 306.65472, 299.20206, 291.8284, 284.4545, 277.0803, 269.70587, 262.48975, 255.11479, 247.97748, 240.36407, 232.59175, 225.21571, 217.68079, 210.38353, 203.36365, 196.1452, 189.00584, 182.02489, 175.12303, 168.3003, 161.15996, 154.33675, 147.67198, 140.92766, 134.34183, 127.83512, 121.64562, 115.059166, 108.393135, 101.56816, 94.90169, 88.15563, 81.48873, 75.05972, 68.90832, 62.63767, 56.446205, 50.333935, 44.459633, 39.06148, 33.504406, 27.867794, 22.151632, 17.467438, 12.624343, 6.907756, 2.6996105, NaN, NaN, 500.33005, 495.6567, 489.6367, 482.0322, 474.58588, 466.74316, 458.97937, 451.37375, 443.53015, 435.60703, 428.00055, 420.3938, 412.7075, 405.25867, 397.80954, 390.59793, 383.3068, 376.17392, 368.96152, 361.98666, 354.6549, 347.52103, 340.30765, 332.77692, 325.3252, 318.03174, 310.73804, 303.3648, 295.91202, 288.45895, 281.0849, 273.86917, 266.65323, 259.5163, 252.37912, 245.1624, 237.86612, 230.56956, 223.59003, 216.21365, 208.48009, 200.94452, 193.56734, 186.03123, 178.65352, 171.35487, 164.29398, 157.23283, 150.40948, 143.42722, 136.36536, 129.46196, 122.71703, 116.13059, 109.46459, 102.95709, 96.92557, 91.0526, 85.17946, 79.306145, 73.43267, 67.55903, 61.447083, 55.176197, 49.063885, 43.18954, 38.029503, 33.107502, 28.502943, 23.580713, 18.896545, 13.974084, 8.495722, 3.6524096, NaN, NaN, 499.0633, 494.54837, 488.92438, 481.08218, 473.4774, 465.79306, 457.95, 449.86896, 442.10455, 434.41907, 426.73328, 418.8095, 411.12314, 403.43652, 395.74957, 387.6661, 379.8201, 371.736, 363.73083, 355.72537, 347.8385, 339.99097, 331.74677, 323.42294, 315.41592, 307.64642, 299.79736, 291.8687, 284.09833, 276.56552, 268.71527, 261.02332, 253.25175, 245.71783, 238.34225, 230.49052, 222.63852, 215.18279, 207.56815, 200.03255, 192.53633, 184.84152, 177.22575, 169.84772, 162.39006, 155.17017, 147.95003, 141.047, 134.14375, 127.55768, 120.81268, 114.384895, 108.11562, 102.08424, 96.13205, 90.10031, 83.98904, 77.718834, 71.13094, 64.46346, 58.11329, 51.60415, 45.094803, 38.744026, 33.26632, 28.106028, 22.945604, 18.261417, 13.656518, 9.369104, 4.128811, 1.4292132, NaN, NaN, 499.4202, 494.9845, 489.20206, 480.3301, 471.14087, 462.5058, 454.26648, 446.10605, 438.183, 430.1012, 422.01907, 413.61966, 405.29916, 396.9783, 388.57788, 380.41486, 372.41003, 364.48416, 356.55798, 348.79004, 341.10107, 333.17398, 325.08804, 316.92252, 308.75668, 300.5112, 291.94827, 283.70212, 275.2971, 266.81238, 258.56525, 250.23846, 242.06996, 233.98044, 226.12856, 218.51431, 210.74115, 203.12633, 195.7492, 188.21317, 180.59752, 172.9816, 165.6034, 158.14558, 151.00487, 143.94327, 136.80206, 129.42256, 122.67761, 115.69438, 108.94899, 101.88593, 94.74326, 87.917816, 81.56836, 75.139336, 68.78948, 62.915688, 56.96235, 50.45317, 44.142242, 37.9502, 32.15491, 26.677025, 21.675348, 16.51476, 11.671627, 7.1459727, 2.8584192, NaN, NaN, 500.21268, 495.46014, 489.36087, 481.0434, 472.6464, 464.32825, 455.85132, 447.69098, 439.37183, 431.1316, 422.89102, 414.88785, 406.72586, 398.72205, 390.63867, 382.555, 374.23325, 366.1489, 358.14352, 349.9793, 341.65622, 333.3328, 325.16757, 317.00204, 308.99475, 300.7493, 292.66208, 284.81244, 277.27963, 269.5087, 261.73746, 254.12453, 246.432, 238.89783, 231.52197, 224.06656, 216.69019, 209.1549, 201.93665, 194.3215, 186.46808, 178.4557, 170.52235, 162.74736, 154.89275, 147.43454, 140.0554, 132.83472, 125.77248, 118.8687, 111.96469, 104.90173, 98.235344, 91.56874, 84.90192, 78.472984, 71.964485, 65.6939, 59.740643, 53.62845, 47.952675, 42.157665, 36.600655, 31.20227, 26.12131, 20.881435, 16.117798, 11.195255, 5.1610093, 1.8262182, NaN, NaN, 502.233, 498.03497, 492.56946, 484.72742, 477.1227, 469.20084, 461.12024, 453.11853, 445.0373, 436.8765, 428.71536, 420.55392, 412.0752, 403.83386, 395.82993, 387.58795, 379.58337, 371.57852, 363.41483, 355.4886, 347.5224, 339.35776, 331.35132, 323.5824, 315.4961, 307.568, 299.56033, 291.71094, 283.62335, 275.53546, 267.52655, 259.27942, 251.26987, 243.0221, 235.17053, 227.23935, 219.14925, 211.93132, 204.71315, 197.33607, 190.15704, 183.01744, 175.79825, 168.3408, 160.64507, 152.55232, 144.69731, 136.76263, 129.14507, 121.60656, 114.14714, 107.00489, 99.94175, 93.11646, 86.449684, 80.0208, 73.98857, 68.35304, 62.71736, 57.081524, 51.286766, 45.015545, 39.61738, 34.13968, 28.741226, 23.34263, 18.182074, 13.735951, 8.495755, 3.4936242, NaN, NaN, 500.96643, 496.60992, 490.74832, 482.74774, 474.82608, 466.82492, 458.90265, 450.90085, 442.5818, 434.50012, 426.3389, 418.2566, 409.85703, 401.53632, 393.2153, 384.89392, 376.81, 368.80502, 360.87897, 352.87338, 344.9071, 337.05942, 329.36996, 321.5217, 313.99023, 306.29993, 298.3715, 290.60132, 282.75156, 274.90152, 266.97186, 259.1212, 251.19093, 243.41898, 235.64673, 228.27075, 220.8152, 213.35938, 206.06192, 198.60556, 191.42657, 183.73169, 176.19518, 168.73773, 161.28001, 153.66335, 146.12573, 138.74654, 131.52577, 124.22541, 117.16286, 110.0207, 103.43382, 96.84673, 90.25943, 83.75128, 77.3223, 70.89312, 64.78124, 58.589806, 52.43787, 46.484207, 40.60976, 35.608406, 30.289371, 24.176281, 19.412708, 14.569629, 8.853059, 3.6921294, NaN, NaN, 498.2344, 493.71942, 487.7785, 480.09467, 472.88586, 465.67682, 458.46753, 451.4164, 444.36508, 437.15503, 430.02396, 422.89264, 415.7611, 408.31232, 400.9425, 393.41394, 386.28137, 378.99005, 371.85696, 364.72363, 357.5108, 350.29773, 343.16364, 336.1086, 329.0533, 321.99777, 315.17984, 308.20312, 301.22617, 294.40756, 287.4301, 280.61105, 273.31598, 266.17923, 259.04224, 251.90501, 244.60892, 237.39188, 230.17458, 223.03633, 215.89784, 208.75911, 201.69946, 194.40158, 187.57942, 180.75702, 173.9344, 166.87355, 160.05048, 153.22716, 146.32428, 139.42117, 132.75589, 125.93167, 119.34529, 112.758705, 106.01318, 99.66426, 93.6326, 87.442024, 81.60842, 75.97309, 70.17885, 64.2257, 58.35175, 52.47763, 46.841496, 40.96705, 36.20386, 31.281782, 25.724453, 20.246368, 15.403302, 10.163134, 3.8112342, NaN, NaN, 501.0864, 496.6507, 490.9475, 482.94693, 475.02527, 467.10327, 459.02255, 450.9415, 442.86014, 434.69925, 426.22107, 417.6633, 409.18442, 400.70517, 392.14633, 383.6664, 375.18613, 366.78476, 358.38306, 350.29807, 342.09387, 333.84967, 325.68445, 317.5189, 309.4323, 301.42468, 293.25818, 285.2499, 277.32065, 269.39105, 261.46118, 253.61029, 245.91772, 238.22485, 230.84895, 223.4728, 216.01704, 208.71967, 201.58067, 194.52077, 187.5796, 180.59854, 173.45857, 166.39769, 159.33658, 152.11653, 144.89622, 137.99306, 130.77225, 123.392494, 116.09182, 108.790886, 101.807144, 94.981895, 88.31515, 81.96567, 75.85411, 69.74236, 63.630436, 57.597706, 51.64418, 45.769863, 39.33968, 33.94134, 29.336763, 25.04965, 20.60366, 16.87213, 11.4732, 5.2801337, 1.9453284, NaN, NaN, 498.55222, 493.40353, 486.9081, 477.95676, 469.08426, 460.3698, 451.655, 442.9398, 433.90732, 425.19138, 416.63358, 408.07538, 399.7546, 391.51273, 383.58752, 375.8998, 368.3703, 360.60275, 352.8349, 345.38385, 337.85324, 330.4016, 322.87045, 315.4976, 307.8073, 300.27533, 292.74307, 285.05197, 277.28125, 269.35168, 261.26318, 253.17436, 245.32315, 237.47165, 229.61983, 221.84705, 214.3119, 206.85582, 199.47879, 192.02216, 184.48593, 176.71143, 168.8573, 161.16153, 153.54483, 145.92784, 138.78667, 131.64523, 124.42421, 117.04421, 109.981384, 102.99767, 95.934364, 89.10891, 82.20386, 75.45732, 69.34556, 63.392365, 57.359623, 50.929794, 44.85699, 38.664932, 32.075737, 26.51842, 21.754885, 16.435472, 10.321949, 4.5258417, 1.9850307, NaN, NaN, 499.0677, 494.4735, 488.61182, 480.69034, 472.7686, 464.8465, 456.84488, 449.00143, 440.9992, 433.15512, 425.39, 417.54535, 409.5419, 401.85513, 394.08884, 386.48074, 378.79312, 371.18448, 363.57553, 356.12485, 348.7928, 341.34155, 333.8108, 326.4383, 319.2241, 312.00964, 304.79495, 297.73856, 290.52335, 283.3079, 275.77502, 268.16254, 260.6291, 253.17468, 245.95792, 238.42366, 230.7305, 223.35431, 215.73991, 207.96658, 200.51025, 192.97432, 185.27946, 177.74298, 170.28555, 162.9072, 155.52858, 148.07034, 140.69118, 133.70851, 126.96366, 119.98052, 113.39393, 106.80713, 100.06139, 93.712265, 87.4423, 80.85467, 74.18745, 67.91689, 61.527077, 55.57365, 49.778816, 43.904434, 37.553562, 31.123102, 25.724537, 20.484615, 15.641539, 9.4485855, 4.128847, 1.3498247, NaN, NaN, 498.31595, 493.80096, 487.93924, 480.3346, 473.04654, 465.83746, 458.4697, 451.2601, 443.81256, 436.444, 429.07516, 421.46835, 413.70276, 406.01614, 398.567, 391.27603, 383.9056, 376.1386, 368.37134, 360.683, 352.95477, 345.1866, 337.57672, 329.6494, 321.88037, 314.03177, 306.18286, 298.49222, 290.88058, 283.1894, 275.81506, 268.2819, 260.74844, 253.76984, 246.791, 239.73262, 232.7533, 225.85307, 218.4767, 211.33801, 204.15942, 196.8616, 189.40486, 181.94785, 174.5699, 167.19168, 159.73387, 152.19643, 145.1348, 138.23161, 131.1695, 124.26584, 117.60003, 111.09271, 104.82327, 98.79173, 92.60128, 86.331276, 79.90234, 73.63195, 67.32168, 61.209656, 55.653114, 49.778893, 44.22204, 38.82381, 32.79033, 26.99484, 21.91373, 16.991285, 11.592339, 6.1932487, 2.779045, NaN, NaN, 500.21762, 495.86108, 490.0786, 482.3156, 474.71075, 467.34326, 459.97552, 452.4491, 445.0016, 437.47458, 429.86807, 422.499, 414.97116, 407.36383, 399.83545, 392.22757, 384.7779, 377.16943, 369.5607, 362.1102, 354.6198, 347.01022, 339.4004, 331.71097, 323.94202, 316.3313, 308.64102, 300.71262, 292.7839, 284.8549, 277.00485, 269.1545, 261.6211, 254.24599, 246.87062, 239.33638, 231.80186, 224.18774, 216.73198, 209.11731, 201.58168, 194.04578, 186.58893, 179.05246, 171.75374, 164.37541, 156.91748, 149.45927, 142.1595, 135.01816, 128.03528, 120.89344, 113.51328, 106.37095, 99.06963, 92.244255, 85.73612, 79.30716, 72.95737, 67.16301, 61.566936, 55.851635, 50.29494, 44.579327, 38.94294, 33.465176, 28.22544, 23.382532, 18.53951, 13.537581, 7.1857486, 2.6599474, NaN, NaN, 499.06958, 494.31696, 488.05917, 479.18704, 469.99765, 461.20398, 452.5684, 443.77396, 435.13763, 426.50095, 418.02237, 409.70193, 401.85666, 394.09033, 386.3237, 378.47754, 370.31403, 362.46722, 354.69943, 347.0106, 339.40073, 331.7906, 324.49725, 316.8073, 308.87918, 300.8715, 292.8635, 284.85516, 276.45007, 268.20322, 259.87674, 251.86713, 243.7779, 235.52974, 227.51918, 219.82559, 212.05238, 204.19955, 196.58441, 188.88966, 181.5516, 174.25296, 167.11273, 159.73424, 152.51414, 145.13513, 137.99388, 130.61433, 122.99646, 115.61637, 108.394745, 101.33158, 94.58564, 87.91884, 81.48994, 75.29895, 69.10778, 63.154552, 57.042393, 51.24758, 45.651062, 40.0147, 34.45757, 29.535416, 24.771927, 19.849539, 14.927033, 9.210425, 3.7318604, NaN, NaN, 500.694, 496.33746, 490.63422, 482.2375, 473.52353, 464.96765, 456.80756, 448.56793, 440.24872, 432.0084, 423.4508, 414.81363, 406.1761, 397.45892, 388.89987, 380.49902, 372.41483, 364.33035, 356.4833, 348.55673, 340.7884, 333.01974, 325.48862, 317.79868, 310.26703, 302.6558, 294.72714, 286.71887, 278.55173, 270.54285, 262.21643, 253.8897, 245.72124, 237.39383, 228.90746, 220.42073, 212.25095, 204.08083, 195.98972, 188.05695, 180.67918, 173.14249, 165.68486, 158.38564, 150.92747, 143.46904, 135.77228, 128.15459, 120.69532, 113.31515, 106.01406, 98.871445, 91.41112, 83.95051, 76.8865, 70.06037, 63.154633, 56.963085, 51.247643, 45.532043, 39.855976, 34.457615, 29.694233, 24.613173, 19.373198, 14.688863, 9.6074295, 5.0816717, 1.9056418, NaN, NaN, 498.9126, 494.3184, 488.37744, 480.4559, 473.24704, 465.8795, 458.51166, 451.1436, 443.696, 436.01047, 428.32462, 420.48004, 412.3974, 404.23523, 396.2312, 388.06836, 379.7467, 371.74176, 363.73648, 355.8894, 348.0817, 340.1548, 332.38608, 324.61713, 316.92712, 309.39542, 301.78415, 294.41046, 286.9572, 279.4244, 272.5257, 265.70605, 258.8862, 252.14542, 245.08717, 238.108, 230.81136, 223.43512, 216.05862, 208.68185, 201.26517, 194.20518, 187.30362, 180.16382, 173.26178, 166.20084, 159.0603, 152.31624, 145.57195, 138.7481, 131.92401, 125.33776, 118.98937, 112.561424, 106.05392, 99.387474, 92.56208, 86.450775, 80.49804, 74.22763, 68.11578, 62.16251, 56.76473, 51.446182, 45.809963, 40.252975, 34.854614, 29.535501, 24.375034, 18.89686, 13.339141, 8.1782675, 5.0022798, 1.9056449, NaN, NaN, 498.47778, 493.80435, 487.62573, 479.38727, 471.4654, 463.86008, 455.85837, 448.17325, 440.17093, 432.406, 424.72003, 416.87527, 409.1095, 401.5019, 393.81476, 386.12732, 378.43964, 370.5931, 362.7463, 355.137, 347.7652, 340.5517, 333.25867, 325.88608, 319.1475, 312.40866, 305.11462, 297.89963, 290.5258, 283.0724, 275.53943, 267.76828, 259.83826, 251.90793, 243.97728, 236.36357, 228.67027, 221.29396, 213.75873, 206.54051, 199.36171, 192.06366, 184.6067, 177.14946, 169.69196, 162.23418, 155.33151, 148.11125, 141.36682, 134.7015, 128.03598, 121.290886, 114.704285, 108.03812, 101.45109, 94.943214, 88.5145, 82.3237, 75.97397, 69.30653, 62.71826, 56.20916, 50.176147, 43.984188, 38.10959, 32.076046, 26.75685, 22.072668, 17.705963, 13.259767, 7.940083, 3.1760702, NaN, NaN, 498.91415, 493.76544, 487.42838, 478.79382, 469.92123, 461.1275, 452.25418, 443.4597, 434.8233, 426.18655, 417.8664, 409.62515, 401.30432, 393.1417, 385.1372, 377.29095, 369.68216, 362.15234, 354.62228, 346.93338, 339.48203, 331.87183, 324.1821, 316.65063, 309.0396, 301.58685, 293.896, 286.20483, 278.59268, 271.13885, 263.44684, 255.75453, 247.98265, 239.7346, 231.48622, 223.23752, 214.82985, 206.65979, 198.64807, 190.71535, 183.09967, 175.56303, 167.7881, 160.40958, 153.11014, 145.96913, 138.98657, 132.00377, 125.4175, 118.910385, 112.561775, 105.89552, 99.22905, 92.9592, 86.84789, 80.89514, 74.7041, 67.71912, 61.21016, 55.018524, 48.58855, 41.92022, 36.124943, 31.044016, 25.883574, 21.67573, 16.594446, 9.92507, 5.1610966, 2.3820608, NaN, NaN, 498.2415, 493.4096, 486.99332, 478.1211, 469.24847, 460.69235, 451.66055, 442.78677, 434.22958, 425.43433, 416.79718, 408.2389, 400.0765, 392.2308, 384.7018, 377.0933, 369.72226, 362.35098, 355.13794, 347.76614, 340.43372, 333.2992, 326.2437, 319.4258, 312.2113, 305.31366, 298.09863, 290.80408, 283.58856, 276.37277, 269.15674, 262.01974, 255.04112, 248.06227, 240.76593, 233.54865, 226.09317, 218.55809, 211.26071, 203.88374, 196.54617, 189.08936, 181.79092, 174.80957, 167.82799, 160.60814, 153.38803, 146.32637, 139.10577, 131.72621, 124.74316, 117.52179, 110.53825, 104.18938, 97.99903, 91.649765, 85.538414, 79.50625, 73.71203, 67.75889, 62.400917, 57.32064, 52.637146, 47.636005, 42.317204, 36.60132, 30.964664, 24.05757, 17.070845, 11.11606, 5.716906, 1.5880456, NaN, NaN, 498.83627, 494.0836, 487.90497, 479.03275, 470.16016, 461.6041, 453.1269, 444.49088, 436.01297, 427.21777, 418.6599, 410.18097, 401.70163, 393.69748, 385.61377, 377.926, 370.1587, 362.54962, 355.09882, 347.64774, 340.19638, 332.824, 325.13428, 317.2857, 309.5954, 302.14267, 294.61038, 287.07782, 279.86215, 272.48764, 265.43005, 258.21362, 251.15555, 243.78001, 236.32489, 228.71086, 220.93793, 213.48198, 205.70847, 198.3313, 190.83485, 183.53648, 176.23784, 168.93893, 161.79846, 154.97511, 148.07217, 141.01033, 134.10693, 127.12395, 120.22008, 112.91919, 105.30059, 97.9198, 90.776855, 83.95113, 77.363304, 70.93401, 64.107635, 57.43979, 51.406788, 45.53238, 39.73719, 34.180008, 29.019629, 23.779726, 17.904524, 13.140724, 8.615011, 4.724406, 1.7071508, NaN, NaN, 500.26294, 495.5895, 489.4109, 481.25168, 473.56747, 465.16998, 456.85138, 448.6909, 439.97543, 431.89352, 423.8905, 415.96643, 408.1213, 400.35513, 392.74716, 385.29742, 377.6889, 370.23862, 362.39175, 354.78238, 347.29163, 339.60245, 331.91296, 323.90607, 316.13672, 308.28778, 300.7557, 293.06476, 285.21497, 277.52344, 270.06952, 262.77396, 255.4781, 248.34062, 241.36151, 234.38217, 227.00601, 219.78822, 212.64949, 205.1139, 198.01434, 190.79553, 183.73514, 176.91249, 169.93095, 162.15578, 154.38031, 146.28716, 138.59044, 131.4489, 124.14839, 116.92698, 109.5466, 101.8485, 94.626305, 87.40386, 80.49864, 73.83132, 67.56066, 61.845463, 56.24918, 50.61305, 45.135536, 39.578487, 34.180065, 28.62272, 23.224012, 18.301535, 13.06135, 6.8682303, 2.3423703, NaN, NaN, 498.28357, 493.29324, 487.03534, 478.3215, 469.2904, 460.41736, 451.38547, 442.43243, 433.39978, 424.44595, 415.80872, 407.40884, 399.1671, 391.5591, 384.1093, 376.65924, 369.6052, 362.47168, 355.3379, 347.88678, 340.47504, 333.18195, 325.4922, 317.64362, 309.71545, 301.5491, 293.54102, 285.37405, 277.44464, 269.7528, 262.0607, 254.44762, 246.91354, 239.22058, 231.68596, 224.07173, 215.98132, 208.44585, 200.51346, 192.73943, 184.76677, 177.07149, 169.05855, 161.28333, 153.34912, 145.732, 137.95589, 130.65561, 123.51377, 116.37169, 109.149994, 102.32486, 95.9757, 89.62634, 83.435524, 77.3239, 71.132706, 65.02071, 58.90853, 52.875553, 46.802704, 40.769367, 34.815243, 29.178514, 23.859203, 18.539755, 13.458363, 8.615042, 4.2480154, 1.3895475, NaN, NaN, 499.90805, 495.39304, 489.45206, 482.24344, 474.95532, 467.27087, 459.5069, 451.58417, 443.42343, 435.0247, 427.101, 418.7016, 410.53958, 402.37723, 394.76932, 387.1611, 379.9489, 372.73645, 365.28598, 358.23154, 351.13724, 344.1616, 337.1064, 329.8132, 322.2819, 314.98813, 307.8527, 300.717, 293.66037, 286.3656, 279.07056, 272.01318, 265.27277, 258.2149, 251.07748, 243.7812, 236.40536, 228.55336, 220.54243, 212.29323, 204.40063, 196.2301, 188.6939, 181.07808, 173.5413, 165.92493, 158.62563, 151.08803, 143.70885, 136.48811, 129.42581, 122.36329, 115.45923, 108.872375, 102.28532, 95.69805, 89.50741, 83.47532, 77.44306, 71.09312, 64.90173, 58.5514, 52.518402, 46.485226, 40.61065, 34.89468, 29.654903, 24.176811, 19.016155, 13.378983, 7.503454, 3.056996, NaN, NaN, 501.53256, 497.17596, 491.39346, 482.759, 474.04495, 465.64743, 457.48724, 449.1683, 440.53207, 431.89548, 423.10004, 414.30423, 405.7458, 397.02847, 388.62784, 380.14758, 371.90475, 363.82013, 355.73517, 347.7292, 339.68326, 331.59735, 323.98682, 316.21744, 308.36847, 300.67776, 292.82822, 284.8198, 276.65244, 268.56406, 260.3961, 251.98984, 243.50397, 234.8591, 226.68977, 218.67876, 210.66742, 202.7351, 194.96114, 187.34554, 180.08665, 172.62918, 165.09209, 157.79274, 150.73119, 143.66937, 137.24213, 130.57661, 123.67282, 116.84815, 110.10262, 103.118774, 96.1347, 89.30911, 82.642044, 76.05413, 69.862885, 63.433323, 57.003555, 50.25605, 43.627407, 37.197018, 30.766426, 24.732601, 19.41316, 13.7759905, 7.9798656, 2.9775982, NaN, NaN, 502.04837, 497.5334, 491.5132, 482.79953, 474.16467, 466.00482, 458.0823, 450.31796, 442.4741, 434.62994, 427.02316, 419.3369, 411.5711, 403.9635, 396.1971, 388.50967, 380.50494, 372.57916, 364.57382, 356.56815, 348.2451, 340.2388, 332.23218, 324.0667, 315.74234, 307.41763, 299.0133, 290.68793, 282.12433, 273.63968, 265.47186, 257.54166, 249.2146, 241.44237, 233.66986, 225.97636, 218.3619, 210.5885, 202.89415, 194.88219, 187.14757, 179.373, 171.99481, 164.85439, 158.11041, 151.52492, 144.85986, 138.11523, 131.29103, 124.06983, 117.24516, 110.49963, 103.912605, 97.72219, 91.61096, 85.737656, 79.62607, 73.75242, 68.11674, 62.322136, 56.328922, 50.613373, 44.81828, 39.419964, 34.418457, 29.416826, 24.494467, 19.492594, 14.649393, 9.647279, 4.803846, 1.7865676, NaN, NaN, 498.48492, 493.96985, 488.108, 480.34476, 472.97736, 465.29276, 457.84558, 450.00198, 441.68268, 433.4423, 425.2808, 417.119, 409.0361, 400.55667, 392.39386, 384.07224, 375.59177, 367.19022, 358.6298, 350.2275, 342.18164, 333.858, 325.53403, 317.28897, 308.80576, 300.32217, 292.0761, 283.90903, 275.7416, 267.41528, 259.1679, 250.92021, 243.22734, 235.37556, 227.68211, 219.90906, 212.21503, 204.1241, 196.11217, 188.41725, 180.8807, 173.50256, 166.28284, 159.22153, 152.0013, 144.54277, 137.32202, 129.9423, 122.8004, 115.89632, 109.071365, 102.246185, 95.500145, 88.75388, 82.08677, 75.26069, 68.355, 61.84599, 55.57491, 49.46241, 43.54819, 37.752888, 32.354374, 27.035109, 21.398127, 15.919785, 10.520695, 5.4390683, 2.183585, NaN, NaN, 497.85202, 493.3369, 487.31662, 479.31567, 471.78976, 464.18436, 456.4202, 448.81424, 441.12872, 432.8883, 424.72678, 416.72342, 408.71976, 400.7158, 392.55298, 384.1521, 376.14716, 368.45895, 360.37415, 352.68536, 345.2341, 337.46548, 329.8551, 322.72012, 315.58493, 308.37015, 300.9173, 293.54346, 286.3279, 279.03284, 271.73752, 264.6798, 257.54257, 250.80164, 244.2984, 237.63632, 231.13266, 224.07358, 216.77629, 209.16147, 201.18938, 193.09799, 185.08562, 177.23161, 169.53596, 161.68137, 153.74712, 146.05058, 138.19508, 130.81538, 123.75286, 116.928154, 110.34131, 103.67489, 97.40508, 91.373184, 85.896706, 80.42008, 74.943306, 69.22826, 63.989323, 58.51211, 53.19352, 47.716022, 42.476536, 37.236916, 32.155945, 27.074848, 22.152414, 17.229862, 12.386592, 7.305004, 3.0173159, NaN, NaN, 499.0804, 494.32767, 488.3074, 480.22726, 472.62216, 464.93756, 457.17343, 449.409, 441.56506, 433.72083, 425.7178, 417.7937, 410.0278, 402.18237, 394.2574, 386.41135, 378.40646, 370.1635, 361.9995, 353.67664, 345.47235, 337.7037, 329.93478, 322.1656, 314.79248, 307.41913, 300.20407, 292.9095, 285.61462, 278.3988, 271.02414, 263.56992, 256.35333, 248.89857, 241.44354, 233.59167, 225.66019, 217.96635, 210.19292, 202.33984, 194.08984, 185.68083, 177.5095, 169.73453, 162.67332, 156.00859, 149.50233, 143.23392, 136.72726, 129.98235, 123.475266, 116.96798, 110.77793, 104.50833, 97.84171, 91.17487, 84.19034, 77.52306, 71.173065, 64.66412, 58.631256, 52.36006, 46.088676, 39.975872, 34.259842, 29.178791, 24.177008, 19.333895, 14.252473, 9.250325, 4.4068594, 1.7865762, NaN, NaN, 500.15048, 495.477, 489.3775, 480.42603, 471.39493, 462.52188, 454.0446, 445.17078, 436.2966, 427.42206, 418.62637, 409.98877, 401.35083, 392.9503, 384.62866, 376.54446, 368.38068, 360.05807, 351.57657, 343.09473, 334.45398, 326.3678, 318.20206, 310.2738, 301.79025, 293.8614, 285.93222, 278.00275, 270.15225, 262.14288, 254.4504, 246.83693, 239.3025, 231.92642, 224.70871, 217.3321, 209.87593, 202.4988, 195.20073, 187.90239, 180.56413, 173.02728, 165.49014, 157.87338, 150.09766, 142.40097, 134.62466, 126.68934, 118.67435, 110.89713, 103.51644, 96.84978, 90.34164, 83.59518, 76.848495, 70.7366, 64.86266, 58.909176, 53.11428, 47.31922, 41.325527, 35.291965, 29.337618, 23.78007, 18.222372, 12.982117, 7.741729, 3.1364279, NaN, NaN, 497.73544, 492.90347, 486.7247, 477.8523, 469.2964, 461.21548, 453.37198, 445.4489, 437.44632, 429.76038, 422.3911, 415.2593, 408.28574, 401.07422, 393.70392, 386.4126, 379.35883, 372.06702, 364.93347, 357.56186, 350.1504, 342.46118, 334.6924, 327.1612, 319.31256, 311.46362, 303.45584, 295.36844, 287.12213, 278.7962, 270.23206, 261.90546, 253.6578, 245.33052, 236.84427, 228.67494, 220.82256, 213.28716, 206.14812, 199.2468, 192.86089, 186.03845, 179.29512, 172.71025, 165.96648, 159.22249, 152.47829, 145.57516, 138.5131, 130.89534, 123.356636, 115.262146, 107.167336, 99.5484, 92.24665, 85.02402, 78.51549, 72.32426, 65.73595, 59.38557, 52.955612, 47.001766, 41.206524, 35.64929, 30.330078, 25.24891, 20.008827, 15.086203, 10.004659, 5.0023904, 2.302703, NaN, NaN, 500.7464, 496.7858, 491.3993, 483.79456, 476.5064, 469.05957, 461.61246, 454.24432, 447.03436, 439.74493, 432.376, 424.84833, 417.3204, 409.31668, 401.15417, 392.9121, 384.82822, 376.10992, 367.7083, 359.30637, 350.8248, 342.18436, 333.78137, 325.37802, 317.05362, 308.8082, 300.5624, 292.55417, 284.54562, 276.53677, 268.6862, 261.15253, 253.69792, 246.32233, 239.02579, 231.57036, 224.2733, 217.05528, 209.67839, 202.61852, 195.51875, 188.14107, 180.60446, 172.98824, 165.37173, 157.51692, 149.6618, 141.56833, 133.39519, 126.01528, 118.55575, 110.93722, 103.318405, 96.175514, 89.270485, 82.68271, 76.09472, 69.5859, 63.394382, 57.202686, 51.090183, 44.818726, 38.705856, 32.83098, 27.511684, 22.351044, 16.793285, 11.314776, 6.0743265, 2.4218118, NaN, NaN, 499.47977, 495.04385, 489.26123, 481.26028, 473.3383, 465.25754, 457.17645, 449.412, 441.568, 433.56522, 425.8791, 417.95496, 410.18903, 402.10577, 394.02222, 385.93835, 377.8542, 369.6904, 361.3678, 353.04483, 344.91974, 336.43756, 327.71722, 318.9965, 310.19614, 301.9504, 293.46646, 285.37863, 277.5284, 269.51926, 261.7477, 253.89656, 246.20374, 238.51062, 230.89653, 223.28217, 215.66751, 208.44919, 201.15129, 194.0118, 186.95139, 179.97006, 172.9885, 165.68935, 158.62796, 151.80437, 144.7425, 137.68039, 131.17351, 124.50771, 118.159134, 111.730995, 105.38202, 99.19158, 92.842224, 86.57203, 80.30165, 73.79295, 67.68094, 61.56874, 55.57543, 49.8598, 44.223392, 38.66622, 33.029507, 27.551422, 21.993797, 16.991806, 11.989692, 6.9874554, 2.9379363, NaN, NaN, 499.16357, 494.56924, 488.54892, 480.1519, 471.4376, 462.6437, 454.08716, 445.37177, 436.81448, 428.49457, 420.3328, 412.24994, 403.3743, 394.65677, 386.17664, 377.29987, 368.58124, 360.10004, 352.01483, 343.77075, 335.44708, 327.20233, 319.19513, 311.1876, 303.4969, 295.2509, 287.32172, 279.31293, 271.70035, 264.16678, 256.87085, 249.73329, 242.59546, 235.53671, 228.23976, 220.78392, 213.16917, 205.79211, 198.57344, 191.3545, 184.29399, 176.99522, 169.77554, 162.71428, 155.4941, 148.74974, 142.0845, 135.3397, 128.1979, 120.57971, 112.961235, 105.263115, 98.12027, 91.61213, 85.26253, 78.753975, 72.40397, 66.371284, 60.100277, 53.749695, 47.75615, 41.881516, 36.40366, 30.131737, 24.097805, 18.619476, 13.299798, 8.059384, 3.2158513, NaN, NaN, 500.82785, 496.5504, 490.847, 482.7669, 475.00336, 467.31876, 459.47543, 451.55255, 443.6294, 436.18134, 428.65375, 421.12592, 413.7563, 406.2279, 398.937, 391.7251, 384.5129, 377.142, 369.92932, 362.63712, 355.30502, 347.69525, 340.08517, 332.55408, 325.02274, 317.6497, 310.4349, 302.90274, 295.05316, 287.20325, 279.67026, 272.37485, 264.9206, 257.9419, 250.88367, 243.74588, 236.3699, 228.67639, 220.50668, 212.25732, 204.16629, 195.9956, 188.14192, 180.28795, 172.67168, 164.49974, 156.16878, 147.91684, 139.74391, 132.04678, 124.50809, 117.60397, 110.85836, 104.5887, 98.63632, 93.001236, 87.28663, 81.730606, 75.777565, 69.348076, 62.918392, 56.567886, 50.05841, 43.31057, 36.403725, 29.337858, 23.065706, 17.269749, 12.108828, 6.788972, 2.6600332, NaN, NaN, 500.82892, 496.23462, 490.21432, 482.6887, 475.4797, 467.71588, 460.03098, 452.42505, 444.81882, 437.2123, 429.60553, 421.91922, 414.3119, 407.02124, 399.6511, 392.04294, 384.51373, 376.98425, 369.296, 361.60745, 354.23566, 346.62582, 338.85715, 331.24673, 323.55676, 316.18362, 308.65167, 300.96085, 293.5076, 286.1334, 278.67963, 271.4635, 264.0092, 256.87183, 249.97215, 242.91364, 235.61693, 228.39926, 221.34, 214.04253, 206.86377, 199.56578, 192.10887, 184.57236, 177.19424, 169.8952, 162.9926, 156.64517, 150.21822, 144.10844, 137.99849, 131.809, 125.61934, 119.27076, 112.68391, 106.33492, 100.303215, 94.112595, 88.00115, 81.81016, 75.46022, 69.34822, 63.077286, 56.964916, 50.931755, 44.819023, 38.150383, 32.037273, 26.400347, 20.525076, 15.284827, 9.965043, 4.9627314, 1.7865971, NaN, NaN, 504.1569, 499.8795, 494.01773, 485.77927, 477.1444, 468.27148, 459.47742, 450.2076, 440.85812, 431.58746, 422.39563, 413.1241, 404.16922, 395.13467, 386.33746, 377.7777, 369.21756, 360.5778, 352.01694, 343.6143, 335.48874, 327.48178, 319.31598, 311.38766, 303.45908, 295.53018, 287.83887, 280.14725, 272.77252, 265.31827, 257.94302, 250.4089, 242.79521, 235.49847, 227.96353, 220.349, 212.4169, 204.2465, 195.75847, 187.19075, 178.82101, 170.33194, 162.00119, 153.98749, 146.2115, 138.59393, 131.21414, 124.23088, 117.32673, 110.97788, 104.708206, 98.43833, 92.247635, 85.6599, 79.2307, 72.32503, 64.942856, 57.71918, 50.81279, 43.82678, 38.15047, 32.91066, 27.194351, 22.19245, 17.349222, 12.18828, 6.5507946, 3.0570636, NaN, NaN, 499.04877, 494.13754, 487.8003, 479.2447, 470.5303, 461.81555, 453.17963, 444.5434, 435.66904, 426.5566, 418.07773, 409.5985, 401.4359, 393.273, 385.10977, 376.94623, 369.0994, 361.25226, 353.3256, 345.3986, 337.43164, 329.2662, 321.259, 313.25146, 305.08508, 297.07693, 288.8306, 280.50464, 271.62323, 262.97937, 254.33513, 245.37328, 236.17311, 227.7657, 219.35794, 211.02916, 202.8587, 194.84657, 187.15146, 178.90071, 171.40335, 163.7867, 156.48715, 148.9493, 141.49051, 133.9521, 126.49278, 119.27126, 112.128845, 104.58936, 97.12897, 89.43019, 82.12799, 74.508026, 66.72902, 59.34663, 52.837204, 46.565735, 40.37346, 34.33978, 29.02047, 24.336185, 19.731192, 14.649698, 9.012269, 3.6922991, NaN, NaN, 500.63388, 495.8811, 489.6231, 481.38446, 473.9377, 466.3322, 458.72647, 451.19965, 443.91028, 436.46216, 429.09305, 421.72363, 414.27472, 406.98404, 399.93085, 392.95667, 385.903, 378.8491, 371.6364, 364.1857, 356.69507, 348.84747, 340.68246, 332.6757, 324.58932, 316.10623, 307.62277, 299.0597, 290.57553, 282.24963, 273.6855, 265.4382, 257.5078, 249.5771, 241.64609, 233.63547, 225.78316, 218.24783, 211.10886, 204.04895, 197.30612, 190.48373, 183.81978, 176.99695, 169.93588, 162.71587, 155.57495, 148.51314, 141.53044, 134.54749, 127.88173, 120.89832, 113.83531, 105.978424, 98.27996, 91.057434, 83.914024, 77.326, 71.05526, 64.546196, 57.759087, 50.217587, 42.913975, 36.165844, 29.496881, 23.939249, 19.810623, 15.602514, 10.679712, 5.836194, 2.3424382, NaN, NaN, 501.42676, 497.2285, 491.8419, 483.9202, 476.3943, 468.47202, 460.62863, 452.70572, 444.62405, 436.54208, 428.45978, 420.53564, 412.69043, 404.84494, 396.9199, 388.83606, 380.5141, 372.58813, 364.82037, 357.21085, 349.6407, 341.87207, 334.42026, 326.73035, 319.35727, 311.90466, 304.1346, 296.9193, 289.86234, 283.04303, 276.54068, 270.19672, 263.61465, 256.87375, 249.57748, 242.20164, 234.74623, 227.1319, 219.51729, 212.14038, 204.5252, 196.75111, 188.81805, 180.488, 171.99895, 163.66823, 155.81323, 148.35468, 141.21324, 134.5477, 128.19934, 122.00952, 115.74014, 109.15312, 102.407166, 95.899086, 89.70828, 83.04105, 75.81798, 68.43589, 61.49013, 54.90137, 49.582577, 45.692623, 42.358322, 37.436153, 31.16419, 26.241755, 21.239803, 15.840735, 10.4415245, 5.121575, 2.0248241, NaN, NaN, 500.79388, 496.43716, 490.65448, 482.49506, 474.573, 466.6506, 458.25256, 450.01263, 441.4554, 433.05634, 425.05313, 417.44583, 409.67975, 401.99265, 393.90897, 385.9835, 377.81995, 369.73532, 361.65036, 353.4066, 345.59845, 337.6711, 329.26782, 321.02274, 312.93588, 304.45227, 295.96832, 287.80118, 279.87164, 272.49686, 265.28046, 258.30167, 251.4813, 244.89862, 238.31573, 231.49469, 224.5941, 217.29668, 209.91966, 202.78036, 195.83916, 188.7787, 181.48, 174.1017, 166.48512, 158.70956, 150.69566, 142.84016, 135.38112, 127.286964, 119.509926, 111.65323, 103.79623, 96.81197, 90.8593, 84.985825, 77.84218, 70.53953, 64.030426, 57.838654, 52.00392, 46.049942, 39.381283, 32.474228, 26.04331, 20.406168, 15.959861, 11.513457, 6.7493467, 2.858574, NaN, NaN, 500.5174, 496.23987, 490.53638, 483.0107, 475.6432, 467.80005, 459.8774, 451.47906, 443.39734, 435.31528, 427.4706, 419.86337, 412.3351, 405.04434, 397.5948, 390.145, 382.8534, 375.48233, 368.34875, 361.29422, 353.84308, 345.91605, 337.4338, 328.47552, 319.59613, 310.79565, 302.23267, 294.06577, 285.81924, 277.57242, 269.64246, 261.63287, 253.7816, 246.32657, 239.42647, 232.68477, 225.62558, 218.32817, 210.79254, 203.33595, 195.83945, 188.30298, 180.84558, 173.62593, 166.32668, 159.10652, 151.56871, 143.95128, 136.57162, 129.66783, 122.7638, 115.62147, 108.16142, 100.93921, 93.87548, 87.76397, 81.01728, 73.952866, 66.33255, 58.950096, 52.242153, 46.685112, 41.445477, 35.88814, 30.092474, 23.899662, 18.580046, 13.816092, 8.496213, 3.335004, NaN, NaN, 498.0227, 493.26984, 487.09097, 478.9314, 471.64294, 463.87888, 455.71838, 447.95374, 440.50574, 433.21594, 425.92587, 418.8733, 412.0582, 405.2429, 398.58588, 391.69086, 384.63712, 377.50385, 370.60815, 363.94998, 357.6087, 351.0294, 344.3706, 338.1873, 332.00375, 325.4236, 318.52615, 311.0735, 303.7791, 296.1673, 288.7931, 281.26004, 273.4888, 266.0345, 258.81784, 251.52159, 244.22511, 236.92836, 229.3934, 222.0168, 214.83824, 207.46114, 199.76643, 192.23012, 184.77286, 177.55333, 170.57156, 163.66891, 156.84537, 150.10095, 143.1976, 136.13533, 128.9141, 121.85132, 115.02638, 108.439316, 101.852036, 95.582016, 90.34362, 85.50196, 79.46957, 73.04011, 66.92797, 61.688847, 56.29082, 49.78125, 42.63636, 36.92027, 32.79188, 29.219172, 23.899687, 17.70668, 11.831091, 6.4317517, 2.7791767, NaN, NaN, 501.7065, 497.2706, 491.32947, 483.17004, 474.69342, 466.05798, 457.42218, 448.9445, 440.22876, 431.51263, 422.71692, 414.0793, 405.44135, 396.96152, 388.5606, 380.00082, 371.91626, 363.75214, 355.66693, 347.8192, 339.89194, 331.8851, 323.87793, 315.94974, 307.70407, 299.29953, 291.1325, 283.12375, 275.4319, 267.73972, 259.88867, 251.958, 244.02702, 235.8578, 227.68826, 219.59772, 211.74483, 203.8123, 196.27612, 188.89833, 181.28227, 173.50725, 165.41457, 157.24222, 148.9902, 140.8172, 132.88194, 125.422516, 117.327934, 110.026665, 102.16958, 93.99471, 86.216385, 79.469635, 73.43706, 67.48368, 62.165188, 56.449635, 50.495766, 44.462337, 38.111164, 31.204042, 25.964003, 22.152979, 17.706696, 13.419116, 8.813838, 4.3672643, 1.6675119, NaN, NaN, 500.4791, 496.04312, 490.18118, 482.0217, 474.41647, 466.81097, 458.80902, 450.8068, 442.80423, 434.56363, 426.56046, 418.6362, 410.87015, 403.34152, 395.8919, 388.52127, 381.0711, 373.69992, 366.48703, 358.9568, 351.14883, 343.4595, 336.087, 328.47638, 320.86548, 313.57144, 305.8807, 298.18967, 290.81552, 283.36185, 275.59067, 268.295, 261.1577, 253.46503, 246.1686, 238.2374, 230.46452, 222.4534, 214.44197, 206.74751, 199.13211, 191.43709, 184.21779, 176.99825, 170.41315, 163.58981, 156.60757, 149.149, 141.61081, 134.23105, 127.24781, 120.18497, 112.96316, 105.66173, 98.518776, 91.216835, 83.597145, 76.45342, 70.18262, 64.943565, 58.950253, 52.67891, 46.169212, 39.7387, 33.863735, 28.941336, 24.336403, 19.25498, 14.173429, 9.329959, 4.565778, 1.7072157, NaN, NaN, 500.24182, 495.72665, 489.7855, 480.83377, 471.72327, 463.16693, 455.40253, 447.63785, 440.03134, 432.3453, 424.97595, 417.76483, 409.9195, 402.39084, 395.02042, 387.5705, 380.35806, 372.98688, 365.69467, 358.1644, 350.4357, 342.7463, 334.9774, 327.446, 319.75577, 311.66885, 303.5023, 295.73187, 288.04047, 280.58667, 272.8154, 264.6473, 256.6375, 248.70671, 241.01353, 233.3994, 225.62634, 218.24959, 210.71393, 203.25732, 195.8401, 188.38295, 181.0842, 173.86453, 166.72395, 159.42442, 152.204, 144.90396, 137.0482, 129.11278, 120.85961, 112.92357, 104.82848, 97.20929, 90.304146, 84.27188, 78.23943, 72.68308, 66.729675, 61.093624, 55.536804, 50.138603, 45.057816, 39.976902, 34.81647, 29.417725, 24.892197, 20.604761, 16.793633, 12.664829, 7.1066933, 3.2159085, NaN, NaN, 500.87592, 496.6776, 490.9741, 482.73544, 474.49643, 466.2571, 458.1759, 449.8567, 441.45792, 432.9003, 424.58008, 416.25952, 407.70087, 398.98337, 390.66174, 382.26056, 373.9383, 365.37787, 356.8964, 348.09747, 339.2585, 330.85522, 322.21375, 313.57193, 305.48474, 297.31793, 289.3887, 282.01422, 274.243, 266.55078, 259.0962, 251.64133, 244.34482, 236.88943, 229.43376, 221.8985, 214.04568, 206.27188, 198.65645, 190.88206, 183.2264, 175.6101, 168.39024, 161.48749, 154.90189, 148.31609, 141.41266, 134.58835, 127.763824, 120.8597, 114.19344, 107.44759, 101.098366, 94.8283, 88.39931, 82.049484, 75.62009, 69.19049, 62.601925, 56.251305, 49.70202, 43.509773, 36.999775, 30.092598, 24.614328, 19.850496, 15.562952, 10.798908, 5.637737, 2.0645413, NaN, NaN, 499.49002, 494.65796, 488.5583, 480.5572, 472.87265, 464.55405, 456.39352, 448.07425, 439.83386, 431.5139, 423.35208, 415.4277, 407.6615, 400.0535, 392.8415, 385.62924, 378.6545, 371.67957, 364.1495, 356.38138, 349.04895, 341.51807, 333.9869, 326.85187, 319.558, 312.50177, 305.2867, 297.83353, 290.14218, 282.45053, 274.75864, 267.14572, 259.29462, 251.3639, 243.35358, 235.6602, 227.88722, 219.95529, 212.34036, 204.8838, 197.58563, 190.52519, 183.54385, 177.19696, 171.0879, 165.13734, 159.26596, 153.23572, 146.49115, 139.90508, 132.922, 125.62127, 118.55836, 111.41584, 104.6699, 98.16184, 91.73294, 85.38322, 78.79517, 72.12754, 65.26123, 58.51377, 51.845474, 44.938797, 38.508232, 32.156857, 26.043472, 20.406296, 14.768962, 9.607886, 5.0819135, 1.8263272, NaN, NaN, 499.21307, 494.8563, 489.23196, 481.3101, 473.3879, 465.3862, 457.46344, 449.22342, 441.22076, 433.2178, 425.21457, 417.36948, 409.3656, 401.44067, 393.75317, 385.98615, 378.1396, 370.5305, 362.7626, 355.15295, 347.3052, 339.21933, 331.2124, 323.04663, 314.88052, 306.87265, 298.9438, 290.69742, 282.4507, 273.8865, 265.16333, 256.5984, 248.27101, 240.02261, 232.01184, 224.31804, 216.38597, 208.21562, 200.12428, 192.27061, 184.41666, 176.32437, 168.07309, 160.37688, 152.68039, 145.22165, 137.92136, 130.70015, 123.55805, 116.0189, 108.6382, 101.17786, 93.95536, 86.33575, 78.636475, 71.57194, 64.983444, 58.950417, 52.9966, 47.280773, 41.247227, 35.53107, 29.735363, 24.495266, 19.334433, 14.41167, 9.568192, 4.4863863, 1.7866257, NaN, NaN, 496.95566, 491.96512, 485.70694, 476.75504, 468.04044, 459.6424, 451.16476, 442.60754, 434.20844, 425.72977, 417.56772, 409.6431, 401.87668, 394.10995, 386.4222, 378.97195, 371.91772, 364.7047, 357.33295, 349.9609, 342.43005, 334.81964, 327.28824, 320.07367, 312.621, 305.6438, 298.74567, 292.00586, 285.26584, 278.5256, 271.78513, 265.04446, 258.54147, 251.80035, 245.13834, 238.39677, 231.73431, 225.15097, 218.48808, 211.9043, 205.20131, 198.29979, 191.39804, 184.25804, 177.5145, 170.85005, 164.10606, 157.20316, 150.30002, 142.99991, 135.54082, 128.0021, 120.22503, 112.606384, 104.987465, 97.923836, 91.41555, 85.224556, 79.27151, 73.318275, 67.44425, 61.966972, 56.648315, 51.805836, 47.122013, 41.96175, 36.404396, 30.60871, 26.24199, 20.525412, 15.443877, 10.52102, 4.4863877, 1.3895997, NaN, NaN, 499.17392, 494.65872, 488.7967, 480.32028, 471.76425, 462.81177, 454.33426, 445.93564, 437.69516, 429.61282, 421.37167, 412.89246, 404.80914, 396.88403, 389.03787, 381.27066, 373.58243, 365.6561, 357.88803, 349.88184, 342.03387, 334.02707, 326.1785, 318.4089, 310.8769, 303.10675, 295.57416, 287.96204, 280.4289, 272.7369, 264.9653, 257.1141, 249.2626, 241.56944, 233.71735, 226.1029, 218.8848, 211.66644, 204.52715, 197.14963, 189.8115, 182.35411, 174.89644, 167.75587, 160.6944, 153.39465, 146.41203, 139.82593, 133.16028, 126.33568, 119.0347, 111.49538, 104.1145, 96.73336, 89.74882, 83.00215, 76.017136, 69.349396, 62.840206, 55.933887, 49.30519, 43.112923, 36.76168, 30.410242, 24.376192, 18.500763, 12.783968, 6.9876094, 2.7791915, NaN, NaN, 497.98593, 493.31226, 487.29178, 478.81528, 470.41763, 462.17813, 453.4629, 444.90576, 436.42752, 428.42438, 420.1832, 412.10016, 403.85834, 395.45764, 387.2944, 379.21008, 371.36325, 363.51608, 355.82718, 348.138, 340.56744, 333.27405, 325.74258, 318.29013, 310.6788, 302.82935, 294.9003, 287.05026, 279.1206, 271.26993, 263.41898, 255.48842, 247.71617, 239.94362, 232.01215, 224.08037, 215.98964, 208.13657, 200.12454, 192.19154, 184.61523, 177.39566, 170.33452, 163.51115, 156.68756, 149.86375, 143.03972, 136.2948, 129.39096, 122.40752, 115.582565, 108.757385, 101.45577, 94.55076, 87.88362, 81.21626, 74.70745, 68.357185, 62.24487, 56.05299, 50.33724, 44.780106, 38.984653, 33.34782, 27.949018, 23.185251, 18.58017, 14.292588, 9.846112, 5.3995395, 2.143952, NaN, NaN, 500.0853, 495.41165, 489.312, 480.67715, 471.9627, 462.77252, 453.34424, 444.47018, 435.83344, 427.5133, 419.03433, 410.7135, 402.23386, 394.46713, 386.70013, 379.0121, 371.16522, 363.39734, 355.78772, 348.25705, 340.4883, 332.63998, 324.79135, 317.02173, 309.09323, 301.1644, 293.2353, 285.14728, 277.13824, 268.89102, 261.03995, 253.02998, 244.9404, 236.69185, 228.20503, 219.79718, 211.07169, 202.82178, 194.80954, 186.797, 178.98247, 171.44534, 163.98727, 156.13222, 148.27686, 139.94508, 132.16844, 124.788315, 117.566635, 110.424065, 103.43998, 97.01123, 90.66166, 84.23251, 77.48566, 70.57983, 63.832527, 57.085007, 50.654804, 44.780125, 38.86558, 33.14935, 27.591751, 22.033998, 16.793695, 12.109068, 7.1861234, 2.6600862, NaN, NaN, 500.28372, 495.37244, 489.19357, 480.24182, 471.3689, 462.65405, 453.8596, 444.98553, 436.19034, 427.23627, 418.51956, 409.88174, 401.00577, 392.12946, 383.56976, 374.77194, 366.3701, 357.88858, 349.72385, 341.55878, 333.15555, 324.9898, 316.98233, 309.13312, 301.28357, 293.43375, 285.74222, 278.209, 270.6755, 263.37964, 255.92491, 248.3906, 240.61807, 233.1625, 225.70668, 218.09193, 210.55624, 203.33757, 196.43597, 189.69281, 182.83041, 175.69011, 168.54956, 161.3294, 154.10901, 146.88837, 139.4294, 131.81145, 124.351944, 117.05088, 109.74956, 102.52734, 95.06677, 87.685295, 80.30355, 72.92155, 66.17432, 59.50625, 52.996735, 46.804565, 40.890076, 35.01511, 29.298767, 24.296835, 19.771173, 15.483611, 11.354762, 6.5111995, 2.8586009, NaN, NaN, 500.2843, 495.68988, 489.59024, 480.87613, 472.39935, 463.76376, 455.44473, 447.12537, 438.88492, 430.8026, 422.64072, 414.71628, 406.71225, 399.02496, 391.2581, 383.41168, 375.7235, 368.03506, 360.42557, 352.57797, 344.7301, 336.88193, 329.11273, 321.42255, 313.8906, 306.517, 298.98453, 291.53107, 284.07733, 276.38544, 268.69327, 261.15942, 253.46667, 245.37708, 237.36649, 229.75217, 222.21689, 214.602, 207.22482, 199.76804, 192.54898, 185.40901, 178.42746, 171.44568, 164.30496, 157.24336, 150.1815, 143.35745, 136.21577, 128.67705, 121.53486, 114.23369, 106.53543, 98.75752, 91.13806, 83.51831, 76.61267, 69.94493, 63.038837, 56.211887, 49.22594, 42.636703, 36.602997, 31.680632, 27.790293, 23.741085, 19.532999, 15.245428, 10.71956, 5.7965727, 2.699794, NaN, NaN, 499.25507, 494.6606, 488.7986, 481.11435, 473.98434, 466.53723, 459.0898, 451.72137, 444.35266, 436.9837, 429.69373, 422.32422, 415.03372, 407.8222, 400.61044, 393.31915, 386.18613, 378.9736, 371.91937, 364.94412, 357.81012, 350.43808, 343.14502, 335.931, 328.95456, 321.97787, 315.08023, 308.10306, 301.12567, 294.14804, 287.1702, 280.1128, 273.29306, 266.5524, 259.6529, 252.75317, 245.61528, 238.63577, 231.5767, 224.83469, 217.97345, 211.23097, 204.32962, 197.34871, 190.60556, 183.86218, 177.19792, 170.45412, 163.55139, 156.96582, 150.38004, 143.8734, 137.6046, 131.25627, 124.90773, 118.71772, 112.28944, 105.781586, 98.956055, 92.28903, 85.859924, 79.50998, 73.318596, 67.28579, 61.332188, 55.775337, 50.456493, 44.978733, 39.65961, 34.8961, 30.370663, 26.083313, 21.87527, 17.428944, 13.061922, 8.933016, 4.4864078, 1.8660399, NaN, NaN, 499.73083, 494.97797, 488.79904, 480.0057, 471.0535, 461.94247, 452.59335, 443.2438, 434.13153, 425.17737, 416.14355, 407.42633, 399.105, 390.46634, 381.8273, 373.10864, 364.70667, 356.54218, 348.5359, 340.5293, 332.68094, 324.75302, 316.82477, 309.0548, 301.5224, 293.5933, 285.74313, 277.8927, 269.96265, 262.1116, 254.33958, 246.56725, 238.71532, 230.9424, 223.32782, 215.87161, 208.17715, 200.7204, 193.10469, 185.56805, 177.87247, 170.4146, 162.95647, 155.33937, 147.48395, 139.86629, 132.40704, 124.39202, 115.97988, 108.12295, 100.10698, 92.646286, 85.42345, 78.200356, 70.73887, 63.59464, 56.608925, 49.384815, 42.63679, 35.888542, 29.656137, 23.780832, 18.302355, 13.3795395, 9.012426, 5.3598614, 2.501286, NaN, NaN, 499.6521, 495.21606, 489.51248, 481.98666, 474.53983, 466.69656, 458.6153, 450.4545, 442.13492, 433.65652, 425.73245, 417.57037, 409.40796, 401.2452, 393.31992, 385.23578, 376.99283, 368.74954, 360.82297, 352.65833, 344.6915, 336.76404, 328.91553, 321.146, 313.45547, 305.76468, 298.07358, 290.54077, 282.7698, 274.99854, 267.227, 259.37582, 251.60368, 244.14848, 236.61371, 229.23729, 221.86061, 214.2457, 206.55116, 199.01501, 191.67691, 184.3782, 177.3966, 170.25609, 162.87729, 155.41887, 148.11888, 141.0567, 133.99426, 127.16966, 120.344826, 113.361046, 106.61512, 99.94834, 93.28134, 86.93162, 80.18482, 73.59656, 67.32561, 61.371998, 55.25944, 48.987926, 42.55744, 36.36493, 30.48981, 25.329096, 20.327045, 15.404275, 10.560787, 5.7171855, 2.4615858, NaN, NaN, 500.04865, 495.45422, 489.43375, 480.2443, 471.2129, 462.10184, 453.38654, 444.4332, 435.7964, 427.39697, 419.07645, 410.91406, 402.83063, 394.82614, 386.90057, 379.13324, 371.28635, 363.35986, 355.5124, 347.9024, 340.52997, 332.84015, 325.38788, 317.7768, 310.08615, 302.3159, 294.3075, 286.37805, 278.28973, 270.1218, 261.95352, 253.70561, 245.616, 237.44675, 229.51514, 221.5832, 213.49232, 205.0045, 196.83363, 188.90045, 181.4033, 173.86623, 166.17017, 158.31514, 150.53917, 142.7629, 134.58955, 126.49525, 118.6387, 110.94058, 103.718376, 96.813385, 90.06691, 83.558334, 76.89079, 70.14366, 63.555073, 56.8075, 50.93296, 44.899475, 38.82612, 33.824394, 28.504965, 23.42359, 18.659687, 13.260464, 7.7816935, 3.2556424, NaN, NaN, 499.89072, 495.29626, 489.1966, 480.40323, 471.92636, 462.89456, 454.02084, 445.22598, 436.03455, 427.0012, 418.52216, 410.122, 401.64227, 393.08292, 384.68173, 376.2802, 367.87836, 359.47617, 351.0736, 343.14636, 335.3377, 327.48914, 319.8781, 312.50467, 304.8138, 297.20197, 289.7484, 282.45316, 275.23697, 268.09985, 260.72455, 253.5076, 246.21107, 238.9143, 231.53795, 224.39929, 217.18108, 209.88327, 202.74387, 195.36621, 187.90897, 180.92747, 174.18375, 167.67784, 161.17172, 154.82408, 148.15886, 141.41406, 134.51033, 127.84445, 120.94027, 113.95649, 106.73438, 99.591385, 92.76562, 86.17775, 79.430916, 72.20759, 65.30153, 58.79216, 52.48105, 46.447605, 40.731544, 35.332897, 30.410477, 26.123112, 21.597462, 16.992311, 12.307656, 6.90826, 2.938024, NaN, NaN, 498.4654, 493.71246, 487.5335, 479.5323, 472.323, 464.87576, 457.42825, 449.5051, 441.81934, 434.21252, 426.84314, 419.55276, 412.10364, 404.97122, 397.68005, 390.54715, 383.57254, 376.3599, 369.46402, 362.48868, 355.5131, 348.69583, 341.87833, 334.98132, 328.00482, 320.79022, 313.41678, 306.0431, 298.90704, 291.9293, 285.1892, 278.4489, 271.47046, 264.65042, 258.14737, 251.32686, 244.42682, 237.60587, 230.94331, 224.35988, 217.81589, 211.31134, 204.64795, 197.905, 191.08249, 184.18044, 177.27814, 169.97891, 162.91745, 156.09378, 149.34924, 142.60448, 135.78015, 129.03494, 122.13079, 115.2264, 108.32179, 101.496315, 94.59123, 88.00342, 81.65351, 75.38279, 69.66753, 63.713966, 57.919, 52.28264, 46.8049, 41.009457, 35.848988, 31.00597, 26.401028, 21.716581, 17.03203, 12.109164, 7.265585, 3.0571353, NaN, NaN, 500.3663, 495.69263, 489.59296, 480.7996, 472.08508, 463.21176, 454.7342, 446.65247, 438.49118, 430.32956, 422.24686, 413.92612, 405.84277, 397.52136, 389.0411, 380.71902, 372.47586, 364.23236, 355.67148, 347.26877, 338.78644, 330.4623, 321.9793, 313.6545, 305.40866, 297.0039, 288.6781, 280.51053, 272.50125, 264.8089, 256.87833, 248.70952, 240.38174, 232.68819, 224.75636, 216.82425, 208.89182, 200.87976, 192.86739, 184.93404, 177.04004, 169.3441, 162.20328, 155.14156, 147.9209, 140.62062, 133.39944, 126.0193, 118.55953, 111.33758, 104.11537, 96.81354, 89.90831, 83.39971, 77.446556, 71.49322, 65.38095, 58.792194, 52.362, 45.693436, 39.5804, 33.784748, 28.30652, 23.463326, 18.540617, 13.617791, 8.139022, 3.454161, NaN, NaN, 500.52426, 496.00906, 489.98862, 481.27448, 472.71844, 464.0036, 455.12994, 446.0974, 436.82678, 427.39725, 417.9673, 409.0124, 400.29486, 391.49768, 382.77942, 374.14005, 365.5003, 356.7809, 348.29898, 339.97525, 331.61157, 323.36642, 315.121, 306.63736, 297.83618, 289.03464, 280.54993, 272.54068, 264.6897, 256.99704, 249.1455, 240.89706, 233.04489, 225.1131, 217.181, 209.40724, 201.87119, 194.41417, 186.87756, 179.02332, 170.7324, 162.63953, 154.70502, 146.6115, 138.91441, 131.2964, 123.75748, 116.21827, 108.75815, 101.45649, 94.71016, 87.725494, 80.58183, 73.834816, 66.92882, 59.784435, 52.877964, 46.130035, 39.85823, 33.983204, 27.949213, 22.470833, 17.309906, 12.387054, 7.543488, 3.4938605, NaN, NaN, 498.583, 493.8301, 487.73038, 478.69928, 469.9055, 461.50745, 453.10907, 444.6311, 436.3905, 428.5458, 420.46304, 412.45923, 404.53436, 396.6092, 388.36667, 380.83716, 373.4659, 365.93588, 358.4848, 350.87494, 343.22516, 335.21835, 327.44907, 319.28305, 311.11673, 303.18796, 295.02103, 286.77444, 278.60684, 270.201, 262.19135, 254.41928, 246.40901, 238.55707, 230.78412, 222.85225, 214.99939, 207.14624, 199.45145, 191.8357, 184.418, 176.96036, 169.74048, 162.52034, 155.37929, 148.63475, 141.96933, 135.4624, 128.87592, 122.209854, 115.54357, 108.797714, 102.131004, 95.860916, 90.06687, 83.87579, 77.92266, 71.81059, 66.01587, 59.90345, 54.108387, 48.392548, 42.358994, 36.08708, 30.529528, 25.368809, 20.684351, 16.237988, 12.029734, 7.3449707, 3.3747492, NaN, NaN, 498.54285, 493.94836, 487.84866, 478.81757, 470.18225, 461.62576, 452.98972, 444.82867, 436.74658, 428.7434, 420.58145, 412.3399, 404.25653, 396.17285, 388.24734, 380.55933, 372.87103, 365.34097, 357.8899, 350.75565, 343.5815, 336.12964, 328.7568, 321.3044, 314.0103, 306.55737, 299.0249, 291.41284, 283.8798, 276.26718, 268.73358, 261.12042, 253.50696, 245.8139, 238.27919, 230.7442, 223.12962, 215.83205, 209.01016, 202.10873, 195.28639, 187.98782, 180.21298, 172.43785, 164.74176, 157.04538, 149.26936, 141.65176, 134.03387, 126.415695, 118.8766, 111.49596, 103.956314, 97.21008, 90.93986, 85.14568, 79.66884, 74.35061, 68.952866, 63.31683, 57.363102, 51.88552, 45.93146, 40.05662, 34.578575, 29.417965, 24.65421, 20.128538, 15.840968, 11.076897, 5.5980763, 2.0248537, NaN, NaN, 500.20554, 495.69034, 489.6699, 481.58957, 473.8258, 465.50717, 457.1882, 449.02737, 440.5493, 432.15005, 423.98825, 415.9846, 408.05988, 400.13483, 392.13025, 384.28387, 376.35794, 368.11465, 360.02954, 352.18195, 344.57187, 336.88223, 329.35086, 321.81924, 314.28732, 306.8344, 299.22266, 291.7692, 283.919, 276.0685, 267.90048, 259.89078, 251.96004, 244.26694, 236.41492, 228.72124, 221.02728, 213.65031, 206.19376, 198.73694, 191.20052, 183.58447, 176.12683, 168.98628, 162.00417, 155.10117, 148.35661, 141.69121, 135.02559, 128.20103, 121.21753, 113.757614, 106.29743, 99.31319, 92.24933, 84.94711, 77.64463, 70.10375, 62.641983, 55.656246, 49.06721, 42.23979, 35.8885, 30.01338, 24.455679, 18.977226, 14.054432, 8.893312, 4.129086, 1.3499026, NaN, NaN, 500.24423, 495.72903, 489.94626, 482.10364, 474.81525, 467.20972, 459.44543, 451.99777, 445.02527, 437.9733, 430.60413, 423.39316, 416.02347, 408.89124, 401.60028, 394.30905, 386.7798, 379.48804, 371.95825, 364.26965, 356.66003, 348.97086, 341.2814, 333.4331, 325.6638, 317.81488, 309.9657, 302.1162, 294.5836, 286.97137, 279.5175, 272.22195, 265.00543, 257.7887, 250.8096, 243.83029, 236.6921, 229.7123, 222.73227, 215.75198, 208.81114, 201.8304, 194.92874, 187.70952, 180.72806, 173.98438, 167.24046, 160.65503, 154.30742, 147.64221, 140.6594, 133.43826, 126.45495, 119.94756, 112.88443, 106.29724, 100.10668, 93.91594, 87.88375, 81.85138, 75.89821, 69.54797, 63.276924, 56.688145, 50.33731, 43.986282, 37.95262, 32.23636, 27.075708, 21.835527, 16.436415, 10.878354, 5.320143, 1.8263334, NaN, NaN, 497.47095, 492.63885, 486.53912, 477.7457, 468.635, 459.7616, 450.88782, 442.17212, 432.9806, 423.4717, 414.20013, 404.76962, 394.8632, 385.19403, 376.07925, 366.80554, 357.45215, 347.93976, 338.50623, 329.23083, 319.95502, 311.0752, 302.43286, 294.10736, 285.9401, 277.7725, 269.84247, 261.75354, 253.58499, 245.49544, 237.56418, 229.63261, 221.70074, 213.92722, 206.1534, 198.37929, 190.2082, 182.35416, 174.81715, 167.67657, 160.69444, 153.95012, 147.36426, 140.77818, 133.95384, 127.04993, 119.987045, 112.685844, 105.7812, 98.63822, 91.57437, 84.51027, 77.44593, 70.30196, 63.71342, 57.4422, 51.647106, 46.090008, 40.13581, 34.73719, 29.41782, 24.09831, 19.016861, 13.776483, 8.377165, 3.8511562, NaN, NaN, 502.42096, 498.3811, 492.91528, 485.152, 477.6261, 469.70377, 461.70193, 453.69977, 445.61807, 437.45682, 429.216, 421.0541, 413.05038, 404.8086, 396.24945, 387.84848, 379.52643, 371.20404, 362.80206, 354.79605, 346.15558, 337.9111, 329.7456, 321.89688, 314.20645, 306.35715, 298.50754, 290.8955, 283.2832, 275.7499, 267.81982, 259.96875, 252.11739, 244.34502, 236.73099, 229.196, 221.34344, 213.64923, 205.79608, 197.94264, 190.28723, 182.75053, 175.13422, 167.35893, 159.6627, 152.1249, 144.50743, 136.49294, 128.63684, 121.01852, 113.79672, 106.89213, 99.987305, 93.32036, 86.57382, 79.827065, 73.63573, 67.682335, 61.80816, 55.854427, 49.463898, 43.19225, 37.39676, 32.474434, 27.393202, 22.470634, 17.389153, 12.228143, 7.225809, 3.0968065, NaN, NaN, 500.24155, 495.8056, 490.41895, 482.89325, 475.68414, 467.99945, 460.31448, 452.6292, 445.0229, 437.4163, 429.65094, 421.9645, 414.59482, 406.9871, 399.3791, 391.85007, 384.16223, 376.39487, 368.86502, 361.41412, 354.04227, 346.82867, 339.45627, 332.00433, 324.71066, 317.41678, 310.51904, 303.85892, 297.04004, 290.3795, 283.79803, 277.13705, 270.71378, 264.4489, 258.18384, 252.0772, 245.97037, 240.022, 233.99414, 228.12473, 221.85855, 215.43355, 208.84969, 202.26561, 195.84, 189.25551, 182.59148, 175.92723, 169.26276, 162.67741, 156.09187, 149.6648, 143.47559, 137.52423, 131.81078, 126.4146, 121.25634, 116.09796, 110.939445, 105.93953, 100.89981, 95.82029, 90.82001, 85.50211, 80.104706, 75.024666, 69.785736, 64.30854, 58.672424, 53.27431, 47.558506, 42.00132, 36.285202, 30.410135, 25.249464, 19.85047, 14.768933, 9.766672, 5.1613073, 2.1439435, NaN, NaN, 501.38907, 497.11157, 491.4873, 483.48633, 475.5643, 467.40427, 459.4816, 451.7963, 443.95227, 436.18716, 428.34256, 420.1014, 411.54294, 402.82562, 394.1872, 384.91437, 375.79962, 366.52594, 357.48965, 348.37372, 339.25735, 330.1406, 320.86487, 311.82657, 302.94647, 294.30383, 285.66086, 277.5726, 269.80124, 262.02957, 254.099, 245.93019, 237.4438, 229.27434, 221.18385, 213.09306, 204.68465, 196.43454, 188.26344, 180.01268, 172.03928, 163.8672, 156.4089, 148.95035, 141.65022, 134.42918, 127.44595, 120.77993, 114.113686, 107.44723, 100.70118, 93.79618, 87.2878, 81.17609, 74.58793, 68.07894, 61.014076, 54.02835, 47.439323, 40.770695, 34.69729, 28.901583, 23.264507, 17.627275, 12.386892, 7.1463757, 2.9379847, NaN, NaN, 500.27908, 495.76392, 489.58514, 481.34647, 473.34512, 465.50192, 457.3415, 449.18076, 441.17816, 433.413, 425.64752, 417.88174, 410.35342, 402.98334, 395.29596, 387.6083, 379.8411, 371.75656, 363.59244, 355.26944, 347.10468, 338.62247, 330.45703, 322.2913, 314.20447, 306.27594, 298.2678, 290.10074, 282.0127, 273.845, 265.7563, 257.66727, 249.65724, 241.6469, 233.55693, 225.70459, 217.77263, 210.07834, 202.38377, 195.00623, 187.66808, 180.29, 173.229, 166.24712, 159.34433, 152.28262, 145.14133, 137.76172, 130.61992, 123.55722, 116.653, 110.542175, 104.3518, 98.08187, 92.129234, 86.097046, 80.38219, 74.74654, 68.8726, 62.601585, 56.092228, 49.74144, 43.54923, 37.912567, 32.593323, 27.750305, 23.224762, 18.699118, 14.093973, 8.615305, 3.4541059, NaN, NaN, 501.2289, 496.71378, 490.69345, 482.21716, 473.2652, 463.8375, 454.33014, 444.82233, 435.23483, 425.4884, 415.97928, 406.4697, 397.19745, 387.84552, 378.81018, 369.93298, 361.05542, 352.65308, 344.2504, 335.60953, 327.20615, 318.961, 310.95337, 302.78683, 294.69928, 286.5321, 278.52322, 270.6726, 262.6631, 254.49466, 246.4052, 238.31543, 230.62192, 222.8488, 215.15471, 207.46034, 199.76567, 192.46738, 185.16881, 177.79065, 170.61058, 163.54927, 156.56706, 149.34657, 142.36388, 135.1429, 128.08037, 121.17631, 113.795845, 105.85957, 98.31983, 90.70044, 83.23952, 76.96895, 71.65073, 66.09423, 60.22005, 54.10755, 48.074253, 42.19956, 36.602562, 31.600864, 26.916622, 21.517702, 15.801042, 9.607814, 3.414399, NaN, NaN, 501.5848, 497.30734, 491.5247, 483.6822, 476.15628, 468.31323, 460.46985, 452.3885, 444.3068, 436.22482, 427.82553, 419.7429, 411.50146, 403.49744, 395.41382, 387.0129, 378.4531, 369.97223, 361.491, 353.2472, 344.8842, 336.4812, 328.3157, 320.0706, 311.5873, 303.5001, 295.41257, 287.40405, 279.39517, 270.59302, 262.1077, 253.93922, 246.167, 238.31517, 230.62167, 222.68993, 215.07515, 207.46011, 200.00343, 192.5465, 185.6446, 178.58382, 172.07817, 165.25493, 158.51082, 151.6078, 144.30779, 137.48364, 130.57991, 123.43787, 116.4543, 109.073685, 102.08963, 95.58154, 88.75577, 82.08852, 75.34167, 68.75336, 62.323593, 56.290546, 50.3764, 44.343, 39.023933, 33.466557, 28.067814, 22.510136, 16.475916, 11.314928, 6.2332134, 2.34244, NaN, NaN, 501.78232, 497.3464, 491.3261, 483.00833, 474.7694, 466.45093, 457.57755, 448.8622, 440.305, 431.58896, 422.3971, 413.44254, 404.09137, 394.8983, 385.86328, 376.66937, 367.31653, 358.28033, 349.16446, 340.9202, 332.63596, 324.1532, 315.90793, 307.9002, 299.57498, 290.93228, 282.5271, 273.40787, 264.05032, 255.08891, 245.96848, 237.48213, 228.75749, 220.5084, 212.02101, 203.85059, 195.67982, 187.11208, 178.70264, 170.76889, 163.0332, 155.09885, 147.16418, 139.38792, 131.92879, 124.23131, 116.37482, 108.9942, 101.53396, 94.54965, 87.644485, 81.05657, 74.46845, 67.48322, 60.577137, 54.06774, 47.875683, 41.842216, 35.411617, 29.29839, 24.137732, 18.579954, 13.419024, 8.257965, 4.0496206, NaN, NaN, 500.07886, 495.6429, 489.781, 481.2255, 472.82806, 463.95496, 455.2399, 446.84143, 438.6803, 430.51886, 422.43634, 414.512, 406.27036, 398.26614, 390.18237, 382.09827, 374.0931, 366.4047, 358.55746, 350.70993, 342.78284, 334.69687, 326.6106, 318.60327, 310.43707, 301.8741, 293.3901, 284.82642, 276.1038, 267.2222, 258.49884, 249.6958, 240.73375, 232.00925, 222.8878, 214.40051, 205.91287, 197.58356, 189.65054, 181.8759, 174.10095, 166.64308, 159.1056, 151.72653, 144.50589, 137.52306, 130.38127, 123.39796, 116.57312, 109.66869, 103.160866, 96.652824, 89.27151, 82.52491, 75.77809, 69.50732, 63.553875, 57.44149, 51.725853, 45.53373, 38.745995, 32.87105, 27.392908, 22.390999, 17.230171, 12.069212, 6.431708, 2.4615417, NaN, NaN, 500.19745, 495.6823, 489.7412, 481.50256, 473.81815, 465.81656, 458.05234, 449.81244, 442.0476, 434.0448, 426.1209, 418.3552, 410.74768, 402.82288, 395.29404, 387.68567, 380.07703, 372.78516, 365.25522, 357.725, 350.2738, 342.42596, 334.6571, 326.88794, 319.19775, 311.34872, 303.658, 295.4119, 287.0069, 278.91876, 270.8303, 262.6622, 254.41449, 246.40437, 238.63187, 230.77977, 223.00668, 215.2333, 207.77693, 200.47894, 193.41869, 186.35818, 179.6941, 173.10916, 166.60335, 160.01799, 153.35306, 146.92596, 140.41931, 133.75375, 127.2467, 120.739426, 114.07323, 107.248085, 100.184616, 93.75585, 87.32689, 80.89773, 74.07148, 67.245, 60.81521, 54.623363, 48.510715, 42.39789, 36.60244, 31.600758, 26.837135, 22.311594, 17.468359, 12.307407, 6.90812, 2.6997528, NaN, NaN, 500.63303, 496.2763, 490.57288, 482.41348, 474.41223, 465.6184, 457.0619, 448.58426, 439.9478, 431.62796, 423.387, 415.06647, 406.7456, 398.4244, 390.02362, 381.86026, 373.69656, 365.61185, 357.6853, 349.59995, 341.4746, 333.0715, 324.8266, 316.42282, 308.57367, 300.64496, 292.71594, 284.7073, 276.53976, 268.60983, 261.07608, 253.70067, 246.48363, 239.66289, 232.60397, 225.62413, 218.4061, 211.26714, 203.7313, 196.67114, 189.49176, 182.27246, 174.89423, 167.27771, 159.6609, 152.04382, 144.10905, 136.25334, 128.63539, 120.93779, 113.319275, 105.70047, 97.922646, 90.70012, 83.715454, 77.04805, 70.301056, 64.03011, 57.52084, 51.170124, 44.819214, 38.547497, 32.59316, 27.035616, 21.716116, 16.634672, 11.553102, 6.3920026, 2.8188581, NaN, NaN, 501.38535, 496.71182, 490.6915, 483.08667, 475.56076, 467.48, 459.31973, 451.23834, 443.07742, 434.8369, 426.91306, 418.90964, 411.06442, 403.13965, 395.21457, 387.28918, 378.88794, 370.96194, 362.79782, 354.47485, 346.50827, 338.0261, 329.54355, 321.13995, 313.05316, 305.04532, 297.19577, 289.10803, 281.33716, 273.64526, 265.8738, 258.02277, 250.72656, 243.35078, 235.7368, 228.51913, 221.38052, 214.47963, 207.5785, 200.35983, 193.06158, 185.8424, 178.2263, 170.68924, 163.15192, 155.69365, 148.07643, 140.53827, 133.47595, 126.492744, 119.5093, 112.208176, 104.98615, 98.16071, 91.33504, 84.58852, 77.92114, 71.01543, 63.871334, 56.806374, 49.62209, 42.874195, 36.7612, 30.489237, 23.026146, 16.118574, 10.560589, 5.161258, 1.9851147, NaN, NaN, 498.65234, 493.97876, 487.72073, 478.76904, 470.21307, 461.736, 453.57547, 445.49387, 437.80814, 430.1221, 422.35654, 414.66995, 407.0623, 399.53363, 391.9254, 384.31696, 376.7082, 368.78207, 361.01422, 353.4046, 345.7947, 337.9467, 329.93982, 321.77408, 313.68732, 305.7588, 297.5921, 289.42508, 281.01987, 273.01077, 264.7635, 256.67447, 248.74376, 240.73343, 232.40552, 224.31523, 216.06598, 207.89572, 199.96312, 192.18887, 184.29533, 176.28249, 168.66603, 161.52534, 154.78113, 148.43344, 142.56165, 136.68968, 131.21432, 125.81817, 120.10445, 114.39056, 108.67651, 103.04168, 97.96226, 93.04144, 88.27926, 83.59633, 78.43705, 72.72201, 66.29239, 59.783188, 53.27378, 46.843555, 39.77801, 33.585533, 28.186813, 23.105534, 17.706535, 11.989795, 6.193492, 2.3821344, NaN, NaN, 500.43445, 495.84012, 489.74057, 481.10587, 472.70844, 463.7561, 455.04108, 446.32565, 437.76837, 429.6069, 421.28665, 413.20377, 405.04135, 396.87857, 388.87402, 381.02765, 373.1017, 365.09622, 356.6941, 348.29163, 339.65097, 331.08923, 322.05148, 313.25116, 304.2919, 295.17365, 285.89642, 276.5395, 267.1821, 257.6657, 248.4661, 239.26607, 229.907, 220.70615, 211.66353, 203.01715, 194.52905, 186.11995, 177.7105, 169.61806, 161.803, 154.42403, 147.20349, 140.22076, 133.15845, 126.17523, 119.19178, 112.04937, 104.82735, 98.081276, 91.73183, 85.144066, 78.238594, 71.571014, 65.141365, 58.711514, 52.678383, 46.96262, 40.84975, 34.57792, 28.583775, 23.264318, 17.944725, 12.148592, 6.2728925, 2.7791533, NaN, NaN, 499.56323, 494.96887, 488.94852, 480.9475, 473.02542, 464.78613, 456.62573, 448.46503, 440.1455, 431.98413, 423.82245, 415.81894, 407.8151, 399.49396, 390.9347, 382.61285, 374.21143, 365.80966, 357.40756, 348.68802, 340.16632, 331.52533, 323.04254, 314.16296, 305.5209, 296.79916, 288.15634, 279.59247, 271.02826, 262.38437, 254.13664, 245.49203, 237.085, 228.59833, 220.50789, 212.6551, 204.88135, 197.42459, 189.80893, 182.35164, 175.01308, 167.6346, 160.25584, 153.0355, 145.73558, 138.27669, 130.81754, 123.9136, 117.168144, 110.5812, 104.07341, 97.56541, 91.37468, 84.94565, 78.59579, 72.08698, 65.33983, 58.671833, 52.083008, 46.04968, 40.33373, 34.697014, 29.139534, 24.058279, 18.500513, 12.466194, 6.193491, 2.461538, NaN, NaN, 502.29623, 497.86038, 491.9193, 483.6808, 475.4419, 467.12347, 458.4878, 450.01022, 441.13614, 432.7371, 424.25845, 415.77948, 407.61716, 399.53375, 391.37076, 383.1282, 374.96457, 366.6421, 358.24002, 349.8376, 341.55374, 333.15063, 324.7472, 316.3434, 307.62213, 299.13834, 290.6542, 282.32834, 274.0814, 266.07205, 258.30032, 250.21104, 242.28008, 234.74536, 227.2897, 219.75446, 212.4569, 205.07974, 197.623, 190.32466, 182.94672, 175.88586, 168.82477, 161.76341, 154.46379, 147.32262, 140.10182, 132.72208, 125.34207, 117.72372, 110.501884, 103.67663, 97.08925, 90.581024, 84.15196, 78.119576, 72.08701, 66.21303, 60.2595, 53.988255, 47.875595, 41.603973, 35.570335, 29.774696, 23.8995, 18.659317, 13.2602, 7.860941, 3.652596, NaN, NaN, 501.62317, 497.26648, 491.40463, 483.64136, 476.27393, 468.58932, 460.74597, 453.0608, 445.61304, 437.61035, 429.2904, 421.44556, 413.6797, 405.83426, 397.90927, 389.82547, 381.89987, 373.65695, 365.25516, 357.01154, 348.80722, 340.64224, 332.47693, 324.46985, 316.62103, 308.8512, 301.08105, 293.38992, 286.09497, 278.64117, 271.2664, 263.97064, 256.75397, 249.45772, 242.24051, 234.86444, 227.4881, 220.27013, 213.13123, 205.83342, 198.6147, 191.3957, 184.17647, 177.03632, 169.81657, 162.59657, 155.45567, 148.15582, 140.69702, 133.23793, 125.937294, 118.16024, 109.98608, 101.73222, 93.47804, 85.302895, 77.76242, 70.38043, 63.474453, 57.04454, 50.93197, 45.057377, 39.658955, 34.260387, 28.385319, 22.589476, 16.15828, 9.488677, 3.9305098, NaN, NaN, 500.51413, 495.9198, 489.82025, 480.94788, 471.59976, 462.33047, 453.06076, 444.10754, 435.15396, 425.88303, 416.69092, 407.57767, 398.62247, 389.66693, 380.79022, 372.0717, 363.35275, 354.47495, 345.676, 337.03525, 328.55267, 320.46616, 312.30005, 304.37146, 296.44257, 288.4341, 280.5046, 272.9713, 265.7549, 258.6176, 251.71796, 244.8974, 238.15591, 231.65216, 225.14821, 218.80267, 212.45695, 206.11104, 199.60626, 193.18062, 186.67545, 180.17006, 173.26778, 166.36526, 159.30385, 152.16283, 144.78351, 137.24522, 129.4686, 121.69168, 113.59702, 105.422676, 97.486115, 89.94609, 82.326416, 75.18272, 68.197525, 61.370857, 54.067657, 47.002357, 40.730705, 35.17339, 29.61592, 24.37588, 19.69149, 14.1336, 7.622737, 3.0967712, NaN, NaN, 497.9792, 493.22635, 487.28516, 479.99707, 473.10483, 465.57858, 457.8936, 450.44598, 443.07736, 435.62924, 428.4978, 421.2869, 414.15497, 406.94354, 399.57336, 392.2029, 384.99072, 377.7783, 370.88263, 363.82822, 356.37723, 349.00525, 341.633, 334.33975, 326.96698, 319.59396, 312.69635, 305.71924, 298.74188, 291.28854, 283.99353, 276.53964, 269.0855, 261.63107, 254.2557, 246.56282, 238.86964, 231.49345, 224.03767, 216.58162, 209.40294, 202.26366, 194.88615, 187.66704, 180.36833, 173.06938, 165.77016, 158.39134, 150.85356, 143.63289, 136.65004, 129.50824, 122.207466, 114.74771, 107.12897, 99.66866, 92.049355, 84.42976, 77.36552, 69.74538, 62.918762, 56.09192, 49.97932, 44.34287, 39.1826, 33.942806, 28.147123, 21.080933, 14.729091, 8.456454, 3.0570683, NaN, NaN, 498.09793, 493.50354, 487.56238, 479.87817, 472.27295, 464.2713, 456.19012, 448.26706, 440.34372, 432.49933, 424.81308, 417.2058, 409.59827, 402.30743, 394.9371, 387.5665, 379.72006, 372.1904, 364.73972, 357.52658, 350.35278, 342.9806, 335.7667, 328.6318, 321.4174, 314.1234, 306.67065, 299.29688, 291.76425, 284.31067, 277.0154, 269.56128, 262.26547, 254.6522, 246.95934, 239.4248, 231.73137, 224.11697, 216.74023, 209.36325, 201.90666, 194.6878, 187.38936, 180.40799, 173.34705, 165.96849, 158.82771, 151.84537, 144.8628, 137.95932, 131.29369, 124.548485, 117.96178, 111.374855, 104.70835, 98.27974, 91.85092, 85.81876, 79.945175, 74.38892, 68.911896, 63.117207, 57.242966, 51.6861, 46.049694, 40.33374, 34.9352, 29.53651, 24.137682, 18.659313, 13.895395, 9.448972, 4.6054354, 1.9057101, NaN, NaN, 499.08798, 494.4144, 488.39404, 479.52158, 470.49033, 461.37943, 452.4266, 444.028, 435.3914, 426.83362, 418.19626, 409.55856, 401.2375, 392.83682, 384.35654, 376.19296, 367.712, 359.15146, 350.5905, 341.94998, 333.46762, 325.30203, 316.97754, 308.6527, 300.40686, 292.31924, 284.5485, 276.53955, 268.6889, 260.75867, 252.51086, 244.57999, 236.49019, 228.16211, 219.67505, 211.50494, 203.09653, 195.08441, 186.99265, 179.13858, 171.60156, 163.7469, 155.97128, 148.43343, 140.97462, 133.67427, 126.45301, 119.46957, 112.485886, 105.26388, 98.27972, 91.454056, 84.62817, 77.80205, 71.37259, 65.181076, 59.465656, 53.6707, 47.954964, 42.318455, 36.761185, 31.283154, 25.804977, 20.406052, 15.4833765, 10.084179, 4.8436437, 1.8263054, NaN, NaN, 501.0285, 496.75104, 491.1268, 482.65057, 473.85712, 465.14252, 456.586, 448.4253, 440.34348, 432.3406, 424.41666, 416.25464, 408.33008, 400.48447, 392.4008, 384.23752, 376.1532, 368.06857, 359.90436, 351.8191, 343.2975, 334.8152, 326.0947, 317.69098, 309.44547, 301.12036, 292.557, 284.3898, 275.82578, 267.57858, 259.4897, 251.24185, 242.83507, 234.34863, 226.09978, 217.92993, 209.36313, 201.03395, 192.70445, 184.1366, 175.72707, 167.31718, 158.9863, 150.81378, 142.56158, 134.30905, 126.373604, 118.675934, 111.37479, 104.15274, 97.00981, 89.946, 82.96132, 76.77015, 70.8963, 65.339806, 59.94193, 54.46452, 48.35188, 42.31844, 36.205437, 30.17164, 24.137669, 18.341711, 12.783791, 7.146317, 2.7791529, NaN, NaN, 501.1471, 496.55276, 490.53247, 481.81857, 472.7874, 463.9143, 455.04083, 446.2462, 437.60965, 428.97275, 421.52414, 413.20355, 404.88263, 396.3236, 387.68497, 378.96674, 370.7237, 362.79736, 354.87076, 346.94382, 338.85803, 331.08905, 323.31976, 315.6295, 307.85962, 300.08945, 292.5569, 285.10333, 277.5702, 270.0368, 262.82034, 255.5243, 248.06941, 241.09012, 234.11058, 227.05148, 220.2301, 213.09122, 205.95209, 198.73337, 191.3954, 183.93817, 176.56001, 169.1816, 161.88223, 154.58263, 146.64798, 139.03043, 131.25388, 123.39768, 115.46182, 107.68439, 100.065384, 92.4461, 85.4615, 78.39729, 71.88849, 65.61761, 59.584682, 53.630962, 47.67707, 41.802395, 36.086334, 30.449503, 24.733124, 19.334173, 14.411477, 8.932853, 3.7716968, NaN, NaN, 499.84003, 495.4041, 489.5422, 482.175, 474.96594, 467.36053, 459.6756, 451.91116, 444.3049, 436.3022, 428.53687, 420.6128, 413.00537, 405.55618, 397.9482, 390.49844, 383.1277, 375.75668, 368.3854, 361.01385, 353.44388, 346.15106, 338.38235, 330.69263, 323.08188, 315.55014, 307.78027, 300.01013, 292.2397, 284.46893, 276.7772, 269.00586, 261.63074, 254.33469, 247.19698, 239.82109, 232.8415, 225.8617, 219.04028, 212.13931, 205.43643, 198.53502, 191.4747, 184.89015, 178.22604, 171.48239, 164.57983, 157.5977, 150.29794, 142.75987, 134.90411, 127.286125, 119.74721, 111.96993, 104.35109, 97.28754, 90.38248, 83.7153, 77.52416, 71.57097, 65.81605, 60.180035, 54.464485, 48.828163, 43.191685, 36.99932, 30.965553, 25.328583, 19.770855, 14.609973, 9.607762, 4.129011, NaN, NaN, 501.3451, 496.83, 490.73047, 482.5711, 474.49066, 465.8553, 457.37805, 449.21735, 441.05637, 432.97427, 424.81262, 416.49216, 408.09213, 399.69174, 390.89474, 382.33514, 373.7752, 365.29416, 356.81277, 348.33102, 340.00748, 331.52505, 323.12155, 314.7177, 306.3135, 297.98828, 289.50412, 281.25748, 273.0898, 264.92184, 256.51562, 248.34697, 240.0987, 231.92941, 223.60115, 215.35188, 207.02295, 198.93167, 190.60208, 182.66882, 175.21127, 167.75346, 160.37473, 153.07506, 145.5371, 138.31625, 130.77774, 122.6041, 114.66821, 106.57329, 98.47805, 90.382484, 83.08033, 76.1748, 69.74529, 63.394966, 56.965065, 50.69373, 44.898525, 39.42072, 34.101547, 29.099815, 23.780376, 18.222605, 12.347084, 6.3125896, 2.1042182, NaN, NaN, 500.43414, 495.91904, 490.374, 482.37305, 474.45105, 466.4495, 458.28915, 450.1285, 442.20526, 434.1232, 425.9616, 417.72043, 409.3997, 401.15787, 392.5987, 383.88068, 375.71707, 367.2361, 358.91333, 350.74875, 342.3064, 333.9826, 325.65848, 317.25476, 309.3264, 301.08054, 292.91367, 284.5086, 276.02386, 267.6181, 259.2913, 251.04346, 243.11253, 235.2606, 227.24976, 219.31792, 211.22713, 203.37398, 195.3619, 187.34949, 179.41609, 171.40306, 163.46907, 155.53476, 147.67949, 140.06198, 132.52353, 125.22288, 118.08068, 110.93824, 103.79555, 97.12881, 90.69997, 84.27092, 77.92104, 71.17409, 64.42691, 57.44136, 50.931885, 44.977913, 39.10316, 33.307632, 27.511936, 22.11306, 16.237652, 10.520874, 5.2009525, 1.7071975, NaN, NaN, 501.42398, 497.06732, 491.28467, 483.0461, 474.88647, 466.25113, 457.53622, 448.7417, 440.26373, 432.1816, 423.86148, 415.46173, 407.1409, 398.26498, 389.38867, 380.43274, 371.55566, 362.75748, 354.03818, 345.08072, 336.4003, 327.91772, 319.5141, 311.03082, 302.86435, 294.93542, 287.08548, 279.15594, 271.46402, 263.8511, 256.3965, 248.78302, 241.08995, 233.39659, 225.70294, 217.53308, 209.28357, 201.03372, 192.3869, 183.97772, 176.00453, 168.30875, 160.77133, 153.313, 145.8544, 138.55423, 131.33315, 124.27052, 116.96958, 109.58901, 102.44628, 95.22393, 88.080696, 80.93721, 73.55534, 66.570114, 59.425877, 52.678318, 46.48624, 40.532146, 34.974834, 29.258583, 24.018547, 18.460787, 13.061676, 8.05943, 3.2952735, NaN, NaN, 499.79984, 495.2847, 489.26437, 480.94653, 472.78677, 464.5475, 455.99097, 447.59253, 439.1938, 430.79468, 422.39523, 414.2332, 405.99155, 397.9081, 389.7451, 381.2647, 372.784, 364.46143, 356.2971, 347.81534, 339.4918, 331.24716, 323.1608, 314.75696, 306.35278, 298.10684, 289.78128, 281.93115, 274.16, 265.9921, 258.45828, 251.0035, 243.38982, 236.17242, 228.71683, 220.62642, 212.69432, 204.3653, 196.1946, 188.26157, 180.44724, 172.67226, 165.05568, 157.51817, 150.5358, 143.3945, 136.09424, 129.26985, 122.60395, 116.01719, 109.27149, 102.76367, 96.335014, 89.82678, 83.79458, 77.60345, 71.41213, 65.37938, 58.94955, 52.83705, 47.041916, 41.484787, 35.9275, 30.37007, 24.73309, 19.413546, 14.0144615, 8.85344, 4.803932, 1.9454075, NaN, NaN, 499.87888, 494.96768, 488.6305, 479.9165, 470.88528, 461.616, 452.4255, 443.4723, 434.43948, 425.7232, 417.4028, 408.76508, 400.2855, 391.48856, 383.0875, 374.76538, 366.5222, 358.3579, 350.0348, 341.55276, 333.0704, 324.5877, 316.3425, 308.25552, 300.16824, 292.23923, 284.3892, 276.69748, 269.32266, 261.94757, 254.25499, 246.64145, 239.18623, 231.81007, 224.03705, 216.58102, 208.96606, 201.19218, 193.49734, 185.88153, 178.26546, 170.64908, 162.7944, 155.2568, 147.87762, 140.81558, 133.83264, 127.1669, 120.262856, 113.596664, 106.93026, 100.025536, 93.35869, 86.69162, 80.02434, 73.51559, 67.24477, 61.211903, 55.25824, 48.82809, 42.913765, 36.88018, 30.846416, 24.733082, 18.698963, 12.823464, 6.788993, 3.2158668, NaN, NaN, 499.08667, 494.4923, 488.55118, 480.07486, 470.64752, 461.29898, 452.4254, 443.63068, 435.07327, 426.4363, 417.8782, 409.31973, 400.84018, 392.51877, 384.11777, 376.03345, 367.94882, 359.78464, 351.6201, 343.37598, 335.29007, 327.3624, 319.35516, 311.50616, 303.4983, 295.4901, 287.4023, 279.31424, 271.2258, 263.13705, 254.9687, 246.40347, 238.07582, 230.0651, 222.13336, 214.20134, 206.42766, 198.65367, 190.87941, 183.2635, 175.568, 167.87218, 160.09674, 152.24167, 144.46564, 136.45125, 128.59526, 120.58027, 113.2792, 106.057236, 98.83502, 91.61255, 84.23108, 77.80184, 71.76929, 65.73656, 59.94179, 53.988094, 48.192993, 42.080177, 36.32444, 30.608232, 24.256706, 17.904984, 12.267663, 6.6301875, 2.1042144, NaN, NaN, 499.4033, 494.72974, 488.7886, 480.94604, 473.1032, 465.0224, 456.7828, 448.93906, 441.095, 433.1714, 425.16827, 417.24405, 409.3988, 401.39474, 393.6281, 386.099, 378.41104, 370.72284, 363.35138, 355.82114, 348.09244, 340.4031, 333.18912, 325.8956, 318.36398, 310.91138, 303.22064, 295.60892, 287.9969, 280.4639, 272.93063, 265.39706, 257.94254, 250.0912, 242.23958, 234.46695, 226.45609, 218.60355, 210.83003, 203.05623, 195.36145, 188.06305, 180.52638, 173.54482, 166.56299, 159.73962, 152.99538, 146.09221, 139.42686, 132.92, 126.65101, 119.90567, 113.39819, 106.89051, 100.144516, 93.557045, 87.36622, 81.01645, 74.90462, 69.18949, 63.752037, 58.35413, 53.03546, 47.875427, 42.556488, 36.99924, 31.600628, 25.963686, 20.326591, 14.848139, 8.813731, 3.2555664, NaN, NaN, 499.16534, 494.57098, 488.3922, 479.99512, 471.20157, 462.16998, 452.97952, 443.78867, 434.8351, 426.11887, 417.48154, 408.6853, 400.04724, 391.40878, 382.61148, 373.89304, 365.25348, 356.6136, 347.89404, 339.57053, 331.24664, 323.0017, 314.83572, 306.74872, 298.81995, 290.8116, 283.12012, 275.11115, 267.33978, 259.48883, 251.47893, 243.54805, 235.77548, 227.76466, 219.99152, 211.6628, 203.4924, 195.55966, 187.78528, 180.0106, 172.43398, 165.45212, 158.62872, 151.96379, 145.21928, 137.9191, 130.3806, 122.92118, 115.54085, 108.71578, 101.811134, 95.54118, 89.58853, 83.39758, 77.20645, 71.41202, 65.61742, 59.902035, 54.027725, 48.073864, 42.199215, 36.16562, 30.211235, 24.733051, 19.254719, 14.093839, 9.17103, 4.40691, 1.7071927, NaN, NaN, 501.26404, 496.74896, 490.88712, 482.807, 474.80582, 466.8835, 458.80246, 450.32495, 441.45093, 432.735, 424.0979, 415.46048, 406.90192, 397.86752, 389.0705, 380.11456, 371.15823, 362.2808, 353.3237, 344.52478, 335.5669, 326.60864, 317.72928, 309.32526, 301.00015, 292.51614, 284.19037, 275.94357, 268.09293, 260.47992, 252.9459, 245.64957, 238.0357, 230.5802, 223.28307, 215.50974, 207.57747, 199.56557, 191.55336, 183.46149, 175.36931, 166.95946, 159.10466, 151.09087, 143.07675, 135.06233, 127.68244, 120.461006, 113.47739, 106.65227, 99.66818, 93.001335, 86.41364, 79.666985, 73.39637, 67.20494, 60.77518, 54.424603, 48.15321, 42.119793, 36.32437, 31.163923, 25.52698, 19.572292, 13.935029, 9.012221, 4.3275037, 1.5483834, NaN, NaN, 498.6893, 493.61966, 487.124, 478.0139, 468.2696, 458.7625, 449.255, 440.064, 430.47638, 421.12604, 411.93378, 403.13736, 394.02353, 385.54337, 376.90433, 368.34418, 359.62515, 351.14355, 342.82016, 334.655, 326.37057, 317.9669, 309.56287, 301.39636, 293.46744, 285.1417, 276.97424, 268.64783, 260.63834, 252.5492, 244.8563, 237.1631, 229.8662, 222.48972, 215.50958, 208.44987, 201.38994, 194.25043, 187.34866, 180.04999, 172.9494, 165.88824, 159.06487, 152.24126, 145.41743, 138.83144, 132.40392, 125.8175, 119.151505, 112.4853, 106.29505, 100.18398, 94.31084, 88.5169, 82.80216, 77.16664, 71.68973, 66.371414, 60.814827, 55.09932, 49.423344, 43.945683, 38.547264, 33.70444, 28.9409, 24.733013, 19.889866, 14.967204, 11.156031, 7.5035896, 3.4540675, NaN, NaN, 499.75842, 495.1641, 488.90613, 480.03378, 470.44803, 461.17874, 452.3844, 443.51047, 434.79462, 425.52374, 416.88638, 408.4864, 399.61057, 390.57584, 381.937, 373.3771, 364.8168, 356.1769, 347.6952, 339.05457, 330.80997, 322.64432, 314.47833, 305.9949, 297.4318, 288.86838, 280.70105, 272.69202, 264.84125, 256.9902, 249.21817, 241.2872, 233.51457, 225.26573, 217.41318, 209.24303, 201.31052, 193.69504, 186.39659, 179.25656, 172.07661, 165.01543, 158.11267, 151.28905, 144.22714, 137.24434, 130.18196, 123.11933, 115.897736, 108.91397, 102.00934, 95.02511, 88.12, 81.37342, 74.86473, 68.35584, 62.00551, 56.13127, 50.177483, 44.382294, 38.66633, 33.18838, 27.789682, 22.787817, 17.706434, 12.863122, 8.257899, 3.3349612, NaN, NaN, 501.8968, 497.2233, 491.12384, 482.7269, 474.09192, 465.21893, 456.1871, 447.2341, 438.043, 429.16846, 420.2143, 411.10123, 401.9878, 393.34946, 384.71075, 376.0717, 366.8774, 358.55466, 350.4694, 342.3045, 334.06006, 325.57742, 317.1737, 308.76968, 299.96884, 291.40552, 283.3176, 275.07077, 266.9822, 258.89334, 250.96277, 243.11119, 235.41794, 227.88304, 220.34785, 212.89172, 205.356, 197.582, 190.12505, 182.42981, 174.6153, 166.91948, 159.14403, 151.36829, 143.43356, 135.49852, 127.959946, 120.50046, 113.8343, 106.92984, 100.18387, 93.834526, 87.32624, 80.897125, 74.467804, 68.11766, 61.687943, 55.019875, 48.748512, 43.112064, 37.991493, 32.98988, 28.226328, 23.70085, 19.413462, 14.887789, 9.171006, 3.6128697, NaN, NaN, 498.80707, 493.97507, 487.79633, 479.47845, 470.92258, 462.4456, 454.28516, 446.12442, 437.96335, 429.485, 421.24402, 413.16122, 405.0781, 396.91537, 388.67313, 380.50977, 372.26685, 364.1821, 356.09705, 348.2495, 340.52057, 332.75168, 325.14108, 316.89594, 308.72974, 300.95966, 293.34787, 285.8944, 278.51993, 271.14523, 263.77023, 255.99847, 248.54364, 241.08853, 233.3159, 225.38434, 217.61111, 209.59962, 201.8258, 194.21036, 186.51527, 179.05792, 171.6003, 163.98372, 156.92227, 149.86057, 142.87798, 136.21255, 129.46756, 123.19848, 117.008575, 110.9772, 105.26311, 99.46948, 93.834435, 88.04049, 82.32575, 76.45211, 70.73705, 64.94246, 59.147694, 53.194004, 47.875225, 43.112022, 38.904434, 34.696762, 30.409607, 25.884182, 22.152615, 17.54761, 12.148505, 5.95524, 2.0645027, NaN, NaN, 499.4799, 494.80637, 488.62762, 479.99292, 471.041, 462.0094, 452.97745, 443.78662, 434.83313, 425.95844, 417.24188, 408.2872, 399.17365, 390.29745, 381.8964, 373.3365, 364.77625, 356.37415, 347.97174, 339.56897, 331.16586, 322.2867, 313.24863, 305.0823, 296.6778, 287.95575, 279.07477, 270.11407, 261.54953, 253.06392, 244.41934, 236.17096, 228.08089, 220.22845, 212.2964, 203.65012, 195.32077, 187.38776, 179.1371, 170.8861, 162.91246, 154.9782, 147.12297, 139.42613, 131.49095, 124.03161, 117.04814, 110.54061, 104.11223, 97.52492, 90.54055, 83.55595, 76.5711, 69.9829, 63.473877, 57.04402, 50.613968, 44.183712, 38.1502, 32.910427, 27.749914, 22.43048, 17.825483, 13.220386, 7.8211718, 2.7394292, NaN, NaN, 499.51907, 494.6871, 488.42917, 479.8737, 471.31784, 462.524, 453.80896, 445.25204, 436.9325, 428.29562, 420.05463, 412.05103, 403.73013, 395.64664, 387.48358, 379.39948, 371.3943, 363.30954, 354.74887, 346.50494, 338.37958, 330.0557, 322.12787, 314.27905, 306.27133, 297.86688, 289.22418, 280.9776, 272.7307, 264.6421, 256.63245, 248.93973, 241.40533, 233.79137, 226.49437, 218.87984, 211.26503, 203.72926, 196.03456, 188.26024, 180.44595, 172.11569, 163.94376, 155.93019, 148.31303, 140.69562, 133.47467, 126.09475, 119.11136, 111.96901, 104.90578, 98.00103, 91.25479, 84.82582, 78.31727, 71.96726, 65.37892, 58.71099, 52.439762, 46.56527, 41.286022, 35.808167, 30.488945, 25.487164, 20.405865, 15.165642, 10.242887, 6.272836, 2.6997254, NaN, NaN, 499.95428, 495.12234, 488.8644, 480.62585, 472.86227, 464.62305, 456.3835, 448.0644, 439.74496, 431.34595, 423.10507, 414.86386, 406.30533, 398.22195, 390.21753, 382.45053, 374.68326, 366.99496, 359.4649, 351.85532, 344.40396, 337.1109, 329.65903, 321.8105, 314.27878, 307.06393, 299.4524, 291.91986, 284.38705, 276.69537, 269.00342, 261.46976, 254.01515, 246.56026, 239.18442, 232.04625, 224.7492, 217.53122, 210.07501, 202.8565, 195.4791, 188.10141, 180.5648, 172.86925, 165.25273, 157.79462, 150.2569, 143.03629, 135.65672, 128.67368, 122.08716, 115.65916, 109.5484, 102.80254, 96.29457, 90.10387, 84.23046, 78.03939, 71.37188, 64.38663, 57.83774, 51.725258, 46.406456, 41.246292, 36.086, 31.004967, 26.638355, 22.271648, 16.952082, 10.838378, 5.439111, 2.183602, NaN, NaN, 499.35965, 494.4485, 488.0321, 479.87274, 472.18835, 463.71146, 455.15497, 446.5189, 437.88245, 429.3249, 420.84622, 412.5257, 403.96707, 395.88364, 387.95834, 380.03278, 371.86914, 363.6259, 355.46158, 347.37622, 339.48874, 331.71985, 323.8714, 316.33975, 308.33215, 300.72067, 292.95032, 285.1797, 277.40875, 269.5582, 261.78668, 253.69765, 246.08414, 238.54967, 231.25285, 223.95578, 216.73778, 209.51952, 202.6183, 195.71686, 188.6962, 181.39761, 174.33678, 166.72034, 158.94492, 151.48659, 144.02798, 136.88652, 129.66545, 122.6822, 115.69871, 108.47689, 101.88974, 95.381744, 89.349754, 83.63508, 77.92024, 72.205246, 66.25196, 59.74283, 53.43195, 47.557503, 42.000435, 36.681385, 31.362198, 25.645903, 20.247032, 14.689222, 9.051862, 4.764188, 1.5880749, NaN, NaN, 499.00256, 494.01218, 487.67502, 479.67407, 472.14813, 463.98813, 456.0655, 447.7464, 439.58542, 431.3449, 423.34177, 415.2591, 407.01758, 399.0135, 391.40536, 383.5592, 375.71274, 367.94522, 360.25668, 352.4886, 344.68057, 337.07047, 329.46005, 321.84933, 314.39694, 306.6271, 299.09488, 291.40375, 283.71237, 276.09998, 268.88382, 261.42947, 253.89558, 246.91656, 239.85799, 232.56123, 225.26422, 217.72899, 210.35213, 202.81636, 195.24065, 187.46631, 179.85036, 172.3928, 164.69695, 157.23885, 150.09784, 142.87724, 135.81511, 128.99078, 122.40429, 115.97632, 109.78622, 103.6753, 97.64357, 91.61166, 85.18271, 78.991684, 72.64172, 66.92658, 61.1716, 55.218, 49.58176, 44.3423, 39.499653, 35.05384, 30.528542, 25.288595, 20.683683, 15.522883, 10.123754, 4.8832846, 1.6277745, NaN, NaN, 497.45743, 492.3878, 485.81293, 477.41583, 468.85992, 460.22443, 451.90552, 443.82394, 435.90054, 427.8976, 420.13208, 412.4455, 404.99637, 397.86395, 390.5728, 383.59845, 376.38605, 369.1734, 361.80197, 354.50955, 346.97906, 339.68613, 332.47217, 325.41656, 318.04355, 310.51175, 302.97964, 295.2887, 287.67673, 280.22308, 272.6106, 264.9978, 257.54333, 250.16792, 242.95085, 235.97147, 228.8332, 221.29813, 213.84207, 206.38576, 198.6912, 190.99632, 183.53918, 175.9231, 168.54474, 161.3248, 154.02527, 146.96352, 140.13956, 132.99797, 126.17356, 119.428276, 112.524055, 105.46087, 99.032364, 92.68303, 86.333496, 80.539375, 74.745094, 69.1094, 63.15603, 57.043728, 51.407547, 46.485683, 41.801865, 37.117943, 32.195736, 27.03523, 21.715805, 16.158049, 10.282542, 4.6450734, 1.6277728, NaN, NaN, 499.5165, 494.44693, 488.03058, 479.47513, 471.07776, 462.44238, 453.72742, 444.77438, 436.05865, 427.5803, 418.86386, 410.14703, 401.35062, 392.47455, 383.5981, 374.80057, 366.24042, 357.7592, 349.2776, 341.03345, 332.59082, 324.02893, 315.6252, 307.37976, 299.21326, 291.205, 283.27573, 275.18756, 267.17834, 259.32745, 251.63489, 244.02133, 236.4868, 228.87268, 221.3376, 213.72292, 206.10796, 198.41338, 190.79785, 183.26137, 176.12129, 168.90163, 161.6817, 154.30284, 146.60632, 138.83017, 130.73631, 122.80085, 115.02379, 107.40517, 100.103714, 93.04011, 86.37311, 80.023384, 73.67347, 67.24397, 61.052418, 55.336967, 49.541973, 43.826206, 38.665997, 33.108707, 27.233692, 21.596695, 16.435926, 12.069022, 6.193403, 2.2232943, NaN, NaN, 499.318, 494.40683, 488.0697, 479.1974, 470.16623, 461.21393, 452.41968, 443.54584, 434.75085, 426.0347, 417.3182, 408.44284, 399.5671, 390.8495, 382.21075, 373.3339, 365.01147, 356.68872, 348.36563, 339.72513, 331.441, 323.11688, 314.4753, 306.07123, 298.14255, 290.13428, 282.12567, 274.27536, 266.58334, 259.04965, 251.51567, 244.06075, 236.52621, 229.15005, 221.93227, 214.31761, 206.782, 199.08746, 191.23398, 183.38019, 175.68477, 167.75105, 160.21373, 152.99352, 145.93173, 138.79036, 131.49004, 124.03074, 116.967964, 109.825584, 102.60359, 95.46072, 88.555695, 81.57107, 74.66558, 67.99799, 62.044605, 56.01166, 50.296078, 44.580334, 38.94382, 33.862885, 28.62304, 22.906693, 17.348978, 12.346907, 7.900518, 3.533435, NaN, NaN, 499.47562, 494.88135, 488.9403, 480.781, 472.7006, 463.98608, 455.192, 446.4767, 437.7611, 429.12436, 420.408, 411.69128, 402.97418, 393.93973, 385.30112, 376.89996, 368.41916, 359.85876, 351.45657, 342.89548, 334.17548, 325.69293, 317.3686, 309.2025, 301.27396, 293.3451, 285.81238, 278.3587, 270.74615, 263.37125, 256.15466, 248.7792, 241.32417, 233.63094, 226.01674, 218.48157, 210.78748, 202.93445, 195.23978, 187.54482, 179.96857, 172.51105, 164.81523, 157.11914, 149.50209, 142.04346, 134.1878, 126.33185, 118.475586, 110.539665, 102.60343, 94.905, 87.60313, 80.380356, 73.31609, 66.330956, 59.90125, 53.630104, 47.914463, 42.51621, 36.998734, 32.076538, 26.519083, 20.564499, 14.689138, 9.76641, 4.6053567, 1.9056776, NaN, NaN, 500.4254, 495.75192, 489.73172, 481.01794, 471.9869, 463.3516, 454.9536, 446.79297, 438.7905, 430.6292, 422.15067, 413.751, 405.74722, 397.74316, 389.58026, 381.49628, 373.09497, 364.6933, 356.29132, 348.12677, 340.1601, 332.15347, 323.98798, 315.90143, 308.05243, 300.44098, 293.06714, 285.69302, 278.08075, 270.4682, 263.0933, 255.63878, 248.10472, 240.8083, 233.19437, 225.8181, 218.28294, 210.50954, 202.73582, 194.96184, 186.94955, 178.61961, 170.68604, 162.91083, 155.294, 147.43887, 139.90083, 132.44186, 124.90327, 117.443756, 110.14269, 102.92074, 95.698524, 88.63479, 81.49145, 74.66535, 68.31529, 62.20317, 56.170254, 50.137154, 44.540504, 38.66584, 32.71162, 26.67783, 21.279026, 16.356462, 11.910175, 5.6375694, 1.9850774, NaN, NaN, 498.16733, 493.25616, 486.8398, 478.36356, 469.9662, 461.48926, 452.85355, 444.21744, 435.34326, 427.1819, 418.94092, 410.62036, 402.458, 394.6123, 386.68704, 378.99927, 371.3112, 363.46432, 355.2208, 347.21478, 338.8517, 330.44867, 322.12454, 314.2758, 306.506, 298.73596, 290.64844, 282.87778, 275.424, 268.04926, 260.67426, 253.06108, 245.52692, 237.91318, 230.37846, 223.16074, 215.7048, 208.48657, 200.95078, 193.0974, 185.32304, 177.94507, 170.56683, 163.02965, 155.3335, 147.79576, 140.33708, 133.2749, 126.371185, 119.46724, 112.483696, 105.65864, 99.38891, 93.67456, 88.436264, 83.0391, 77.80053, 72.0062, 65.497314, 58.829453, 52.39953, 46.366325, 40.96805, 36.045963, 30.806196, 25.72508, 20.96142, 16.038857, 11.27497, 5.7963653, 2.1438801, NaN, NaN, 499.27576, 494.36462, 488.10675, 479.789, 471.62936, 463.15253, 454.59607, 446.11853, 437.71985, 429.08313, 420.68378, 412.2841, 403.88403, 395.24588, 386.7659, 378.3648, 369.88412, 361.08603, 352.4461, 343.96436, 335.72006, 327.7133, 319.86475, 311.85736, 303.84964, 295.8416, 287.754, 279.66605, 271.4985, 263.172, 255.00378, 247.07317, 239.22156, 231.21101, 223.75539, 216.53745, 208.76398, 201.06956, 193.29552, 185.8385, 178.38123, 171.003, 163.86255, 156.48381, 149.2635, 141.88425, 134.66342, 127.28363, 120.30036, 113.158134, 105.936295, 98.79357, 91.6506, 85.2217, 78.79261, 72.60145, 66.251335, 60.139168, 53.709286, 46.961666, 40.332905, 33.981792, 28.027447, 22.549295, 17.229792, 11.671953, 5.3993535, 1.9056704, NaN, NaN, 499.592, 494.7601, 488.58145, 480.0261, 471.2327, 462.2805, 453.16943, 444.2957, 435.9762, 427.41864, 419.25696, 410.6987, 402.4571, 394.21518, 386.1314, 378.1266, 370.12146, 361.87823, 354.1103, 346.57986, 339.04913, 331.5974, 324.14542, 316.77246, 309.55777, 302.10498, 294.9691, 287.59506, 280.2208, 272.68765, 265.07492, 257.6205, 250.32446, 242.86954, 235.57295, 228.1175, 220.74107, 213.36438, 205.82878, 198.29291, 190.47911, 182.46667, 174.1366, 166.04419, 157.95146, 150.1758, 142.39984, 134.70293, 126.926384, 119.546326, 112.483444, 105.6584, 98.67441, 91.84891, 85.10255, 78.75283, 72.641045, 66.529076, 60.337543, 54.14583, 47.834843, 41.56336, 35.60924, 29.813734, 24.494425, 19.49256, 14.887561, 9.567863, 4.1686263, 0.59552324, NaN, NaN, 499.35373, 494.28418, 487.70944, 478.8372, 469.8853, 460.53693, 451.02966, 441.52197, 432.25156, 422.9807, 413.78867, 404.04153, 394.69016, 385.17987, 376.0654, 366.6335, 357.5975, 348.3233, 338.89014, 330.01147, 321.25134, 312.4512, 303.9678, 295.80124, 287.71362, 279.54642, 271.45816, 263.0524, 255.0428, 247.19151, 239.49855, 231.8053, 224.03244, 216.10065, 208.08922, 200.39479, 192.54141, 184.52908, 176.43709, 168.5828, 160.80754, 153.032, 145.3355, 137.87677, 130.1797, 122.64106, 115.34022, 108.2772, 102.007576, 95.97585, 90.3408, 84.62621, 78.8321, 72.56158, 66.449615, 60.496227, 54.70143, 48.90647, 43.508278, 37.871777, 32.51299, 26.876186, 22.11257, 17.42824, 12.743802, 7.0270543, 2.739389, NaN, NaN, 499.98676, 495.39252, 489.29312, 480.97546, 472.57825, 464.02222, 455.22818, 446.35452, 437.79745, 429.0815, 420.20676, 411.41083, 402.6938, 393.89716, 385.2586, 376.54047, 368.05975, 359.2616, 350.78015, 342.37766, 334.45044, 326.44363, 318.59506, 310.98407, 303.2142, 295.60263, 287.8322, 279.98218, 271.97327, 264.04333, 256.03378, 248.26184, 240.80685, 233.82747, 227.00648, 220.50255, 213.6811, 206.62149, 199.32364, 191.78755, 184.44951, 177.30954, 170.328, 163.58424, 156.99895, 150.1754, 143.1136, 135.97218, 128.9099, 121.76799, 114.38777, 107.00728, 99.15034, 91.68993, 84.78485, 78.27639, 72.085236, 65.89388, 59.86111, 54.38383, 49.660553, 45.215015, 40.13428, 34.656475, 29.019741, 23.62103, 18.777948, 14.172946, 9.012043, 3.5334032, NaN, NaN, 500.22388, 495.23358, 488.73813, 479.78668, 470.99335, 461.64502, 452.21707, 442.78867, 433.59756, 424.80222, 416.00653, 407.36893, 398.81024, 390.09268, 381.61252, 373.132, 364.73038, 356.48697, 348.24323, 340.23697, 332.27005, 323.62894, 315.06677, 306.42496, 298.1792, 290.01242, 282.0832, 273.99506, 265.8273, 257.26273, 248.38055, 239.498, 231.01163, 222.68353, 214.75171, 206.89891, 199.04579, 191.19238, 183.81467, 176.43668, 169.49478, 162.35431, 155.37227, 148.46933, 141.64551, 134.90082, 128.23526, 121.56948, 114.74477, 108.078545, 101.6502, 95.14229, 89.03101, 83.55452, 78.07788, 72.12485, 65.77475, 59.6626, 53.550266, 47.358364, 41.245663, 35.529724, 29.972408, 24.891302, 20.048256, 14.8875065, 9.567828, 4.406815, 1.6277535, NaN, NaN, 499.23322, 494.55975, 488.61877, 480.85562, 473.80515, 466.2791, 458.83203, 451.4639, 444.25397, 436.5684, 428.72406, 420.8794, 412.95523, 405.26846, 397.42294, 389.49786, 381.81024, 373.726, 365.56226, 357.31888, 349.2337, 341.2275, 333.1417, 324.7385, 316.41418, 308.56528, 300.39893, 292.3908, 284.62027, 276.53223, 268.6025, 260.67245, 252.98003, 245.04938, 237.27704, 229.50441, 221.89012, 214.11693, 206.34341, 198.56963, 191.03352, 183.33847, 176.03981, 169.05824, 161.91776, 154.69768, 147.39801, 139.93938, 132.55981, 125.57677, 118.83156, 112.165474, 105.81663, 99.46758, 93.27708, 87.5626, 81.68922, 75.81567, 69.783195, 64.226814, 58.789356, 53.39144, 47.914, 41.9601, 36.482353, 30.925068, 25.129456, 19.651258, 14.093518, 9.250221, 4.4862113, 1.9453603, NaN, NaN, 501.094, 496.579, 490.40042, 481.9244, 473.52725, 464.49597, 455.4643, 446.353, 437.479, 428.44617, 419.33365, 410.0623, 401.1867, 392.70703, 384.06848, 375.4296, 366.55252, 357.27878, 348.32166, 339.20563, 330.00992, 320.97235, 312.09296, 303.0546, 294.49158, 286.16608, 277.84024, 269.27618, 261.18756, 253.25725, 245.40593, 237.63362, 229.86102, 222.00882, 214.31494, 206.54146, 198.60902, 190.75562, 182.74324, 174.49255, 166.43988, 158.10919, 149.77817, 141.28812, 133.2738, 125.89402, 118.8314, 111.92725, 105.102234, 98.594444, 91.92772, 85.498886, 78.9111, 72.95811, 67.08431, 61.607246, 56.130035, 50.25576, 43.984386, 38.18915, 32.949482, 27.947853, 23.025497, 17.467855, 11.274878, 4.6053066, 0.9528306, NaN, NaN, 498.3606, 493.37027, 486.95398, 478.87393, 471.26886, 463.42587, 455.18643, 447.10513, 439.0235, 431.10004, 422.93854, 414.856, 406.6146, 398.2144, 389.49683, 380.7789, 372.0606, 362.94565, 354.06808, 345.58646, 336.94595, 328.1465, 319.90167, 311.81506, 303.72815, 295.87875, 288.34622, 280.97205, 273.59756, 266.14352, 258.76852, 251.23465, 243.7798, 236.404, 229.02794, 221.49297, 213.79909, 205.78763, 197.77585, 189.44644, 181.4737, 173.46097, 165.84464, 158.228, 150.84912, 143.70802, 136.72537, 129.74248, 122.838715, 116.252144, 109.82407, 103.633896, 97.20544, 90.61804, 84.03043, 77.60136, 71.013336, 64.50447, 58.551064, 53.073776, 47.516956, 41.801216, 36.482258, 31.639502, 26.717241, 22.033043, 17.34874, 12.743726, 7.424011, 2.977577, NaN, NaN, 498.83536, 493.84506, 487.66644, 479.42798, 471.34763, 462.87085, 454.23526, 445.837, 437.35916, 428.80176, 420.244, 411.6066, 402.6519, 394.17227, 385.69232, 377.13275, 368.4143, 360.01257, 351.769, 343.68365, 335.91507, 327.74982, 319.6635, 311.73547, 303.80713, 296.03705, 288.66312, 280.89246, 272.96292, 265.42957, 258.05453, 250.44135, 242.43132, 234.26236, 226.01376, 217.92346, 210.15013, 202.21786, 194.68192, 187.14569, 179.68854, 172.07243, 164.21802, 156.12529, 148.11159, 140.49431, 132.9561, 125.65568, 118.593056, 111.76828, 105.57816, 99.62595, 93.51485, 87.32418, 81.92704, 76.13289, 70.2592, 64.70285, 59.46387, 54.14538, 48.70767, 42.674423, 36.402832, 30.607395, 25.28815, 20.206951, 15.205024, 9.726582, 4.3273935, 1.5483439, NaN, NaN, 501.25092, 496.5775, 490.399, 481.68533, 472.33755, 462.8309, 453.4823, 444.45016, 435.3384, 426.54318, 417.82684, 409.34787, 400.86853, 391.9926, 383.51257, 375.0322, 366.3929, 357.7533, 349.1926, 340.31442, 331.8719, 323.31012, 314.90652, 306.18546, 297.30545, 288.58362, 279.94073, 271.1389, 262.416, 254.0892, 246.00002, 238.30707, 230.53452, 222.52371, 214.75056, 206.8978, 198.41013, 190.1601, 182.06839, 174.0557, 166.51872, 159.29884, 152.2374, 145.41373, 138.11375, 130.73416, 122.719475, 115.101265, 108.038284, 101.37189, 94.70527, 88.117805, 81.53013, 74.86286, 68.59226, 62.242092, 56.44739, 50.652527, 44.698723, 38.903526, 32.869995, 27.153852, 21.675734, 16.118073, 10.639658, 5.2404976, 1.7468475, NaN, NaN, 500.4583, 495.7849, 489.76477, 482.08093, 474.55524, 466.55392, 458.39386, 449.9958, 441.59738, 433.43634, 425.1957, 416.63782, 408.3965, 400.31342, 392.38846, 384.701, 377.01324, 369.3252, 361.9539, 354.58234, 346.97275, 339.52136, 331.9112, 324.4593, 317.0864, 309.23755, 301.3091, 293.45966, 285.60992, 277.99774, 270.4646, 262.85187, 255.47676, 247.94278, 240.17061, 232.2395, 224.3081, 216.37639, 208.36505, 200.59137, 192.89673, 185.43977, 177.98257, 170.44576, 162.82932, 155.29193, 147.99232, 140.53375, 133.31296, 126.25061, 119.505455, 112.60136, 105.61767, 98.47501, 91.17337, 83.7921, 77.124916, 70.37814, 64.504295, 58.868427, 53.549923, 48.231285, 42.833122, 37.831757, 33.068436, 28.225613, 23.303284, 18.222044, 13.061281, 7.344592, 2.977569, NaN, NaN, 498.319, 493.64554, 487.70456, 480.17908, 472.4949, 464.57275, 456.6503, 448.72754, 440.96292, 433.1188, 425.43286, 417.6674, 410.13934, 402.69028, 395.08246, 387.7121, 380.3415, 372.9706, 365.59946, 357.91098, 350.61856, 343.24664, 335.71588, 328.50195, 321.1292, 313.67694, 306.22437, 299.00943, 291.7942, 284.42014, 277.04584, 269.59195, 262.2171, 254.9213, 247.38731, 239.93236, 232.31851, 224.46643, 216.61406, 208.76137, 201.06705, 193.53108, 186.07417, 178.93433, 171.79424, 164.8919, 158.06868, 151.0072, 144.50092, 137.91505, 131.40836, 125.139496, 118.94981, 112.998, 106.807945, 100.6177, 94.42727, 88.07791, 81.8871, 75.93423, 70.02086, 64.067635, 58.35238, 52.636963, 47.15954, 41.68197, 35.966087, 30.408827, 24.613237, 19.055668, 13.815536, 8.57527, 3.6524737, NaN, NaN, 498.87283, 494.041, 487.70395, 478.8318, 469.7216, 460.61096, 451.3415, 442.30933, 433.51443, 424.40222, 415.52734, 406.57285, 397.93494, 389.2174, 380.57877, 372.0983, 363.5382, 355.45334, 347.36816, 339.44122, 331.51398, 323.42786, 315.5, 307.88895, 300.51547, 292.98315, 285.4506, 278.3142, 270.93967, 263.72348, 256.34845, 249.13173, 241.51823, 233.82513, 226.68697, 219.70717, 212.48918, 205.35027, 197.97311, 190.35773, 182.74205, 174.88808, 167.27184, 159.73463, 152.35585, 144.9768, 137.59749, 130.29726, 123.39355, 116.4896, 109.58542, 102.76037, 95.69699, 89.34769, 83.31567, 77.28346, 71.33046, 65.37728, 59.26517, 53.073498, 47.15948, 41.443756, 35.96604, 30.805738, 25.724699, 20.405352, 15.16526, 9.925035, 4.684677, 1.7468412, NaN, NaN, 500.10013, 495.2683, 489.01056, 479.98, 471.02832, 462.0762, 453.20297, 444.40854, 435.9307, 427.611, 419.29092, 410.81204, 402.25357, 393.9325, 385.53183, 377.21005, 368.72946, 360.08997, 351.76718, 343.20627, 334.36752, 325.96442, 317.32315, 308.76077, 300.11877, 291.08, 282.19934, 273.23904, 264.43695, 255.63448, 246.91095, 238.34566, 229.46275, 221.13469, 213.04424, 204.95348, 197.10036, 189.40561, 181.55191, 173.6979, 165.68494, 157.67165, 149.49934, 141.16803, 132.91574, 124.58375, 116.64821, 108.95045, 101.56984, 94.82389, 88.395195, 82.12504, 75.93406, 70.13977, 64.504074, 58.86822, 53.152832, 47.754818, 42.197887, 37.117134, 32.115646, 26.87586, 21.238972, 15.998906, 10.520514, 5.3595743, 2.1835473, NaN, NaN, 500.575, 495.90164, 489.88153, 481.48477, 473.1669, 464.61102, 455.89633, 447.18127, 438.6243, 429.82928, 420.95465, 412.15887, 403.3627, 394.80392, 385.7693, 376.73425, 367.77805, 359.05927, 350.49866, 342.01697, 333.33673, 324.8543, 316.37155, 308.44342, 300.83212, 292.9827, 285.21225, 277.5208, 269.51187, 261.34402, 253.17587, 245.48323, 237.7903, 230.09708, 222.4829, 214.70978, 206.93637, 198.9247, 190.99203, 183.1384, 175.6018, 167.9856, 160.28976, 152.5143, 144.73853, 137.04182, 129.66223, 122.52045, 116.17198, 110.140755, 103.63319, 97.204765, 90.696785, 84.10922, 77.36271, 70.77472, 64.26589, 58.233143, 52.279594, 46.405254, 40.570442, 34.854546, 29.694223, 24.216202, 18.896824, 13.736099, 7.9400544, 3.017257, NaN, NaN, 499.06946, 494.2376, 487.8214, 478.87006, 469.36377, 459.93628, 451.14218, 442.5854, 434.02826, 425.3915, 416.59595, 407.95847, 399.47916, 391.39572, 383.23273, 375.22794, 367.30206, 358.97958, 350.73605, 342.1751, 333.81198, 325.3296, 316.76758, 308.2845, 299.95963, 291.55515, 283.3089, 274.98303, 266.5775, 258.33026, 250.00339, 241.8348, 234.22104, 226.60701, 219.15134, 211.93335, 204.55646, 196.70335, 189.2466, 181.94823, 174.72893, 167.58871, 160.36891, 153.30754, 145.92854, 138.31125, 131.01106, 123.86932, 116.965416, 110.29935, 103.633064, 97.12529, 91.014145, 85.22029, 79.66439, 73.87022, 67.996506, 62.122627, 56.248577, 50.453743, 44.777824, 39.220825, 33.425507, 27.709417, 22.548923, 17.467691, 12.54513, 7.1460543, 3.0966542, NaN, NaN, 498.94986, 494.19724, 488.1771, 480.09714, 472.17532, 463.93634, 455.53854, 447.3781, 439.45502, 431.05624, 422.81558, 414.81235, 406.6503, 398.4879, 390.4837, 382.16217, 374.15735, 366.15222, 357.90897, 349.74466, 341.6593, 333.49435, 325.1705, 317.0842, 308.99756, 301.22772, 293.37833, 285.6079, 277.83722, 270.7006, 263.56372, 256.5852, 249.44786, 242.31026, 235.41034, 228.19293, 221.45117, 214.47122, 207.25308, 199.95537, 192.73671, 184.88316, 177.26732, 169.6512, 162.11412, 154.89413, 147.91194, 141.0882, 133.78812, 126.963905, 120.377525, 114.029015, 107.36286, 100.775856, 94.268005, 88.077415, 82.04538, 76.33066, 70.695145, 65.05949, 59.542736, 53.986145, 48.429405, 42.872513, 37.236084, 31.917059, 26.677286, 21.357986, 16.435526, 11.512946, 5.716854, 2.1438391, NaN, NaN, 498.3551, 493.28564, 486.711, 477.83884, 468.6494, 459.61804, 450.03165, 440.99945, 432.2046, 423.1716, 413.97974, 405.10446, 396.30804, 387.5905, 378.79333, 370.47137, 362.3868, 354.6983, 346.61313, 338.28986, 330.28333, 322.5143, 314.50717, 306.6583, 298.8091, 290.72177, 283.03055, 274.94257, 267.2508, 259.8759, 252.42145, 244.88742, 236.87726, 229.34267, 222.04575, 214.9072, 207.7684, 200.86732, 193.64871, 186.42986, 178.8934, 171.35669, 163.42299, 155.489, 147.71338, 139.77878, 132.16125, 125.1783, 118.353806, 111.52908, 104.70414, 98.19642, 92.00596, 85.89468, 79.86259, 73.90969, 68.11537, 62.479645, 56.92314, 51.04896, 45.253998, 39.776413, 34.854404, 29.852882, 25.327593, 20.484629, 15.323965, 10.083775, 4.9228497, 1.6674302, NaN, NaN, 499.78046, 494.94864, 488.53247, 480.61102, 472.68924, 463.9749, 455.49792, 447.09982, 438.5429, 430.1441, 421.9034, 413.74167, 405.4211, 397.57568, 389.49222, 381.40845, 373.32434, 365.63623, 358.02707, 350.25912, 342.49088, 334.56378, 326.08148, 317.28168, 308.32297, 299.83957, 291.35583, 283.1096, 275.02164, 267.09195, 259.16196, 251.46959, 243.93553, 236.16327, 228.54933, 220.93513, 213.24132, 205.4679, 197.61485, 189.92017, 181.82854, 173.89525, 166.51703, 158.97986, 151.68044, 144.61879, 137.7156, 130.89154, 123.511765, 116.52851, 109.54501, 102.95809, 96.52969, 89.86298, 83.434166, 77.00515, 70.73468, 64.543396, 58.51068, 52.239643, 46.32564, 40.768707, 35.21162, 30.130722, 25.129091, 20.127338, 15.046067, 9.567679, 4.2479463, 1.5483271, NaN, NaN, 502.15625, 497.79977, 492.0174, 484.09604, 476.016, 467.46027, 458.74576, 449.8724, 440.8402, 431.41147, 421.98227, 412.6319, 402.80563, 393.1374, 383.70645, 374.51285, 365.3981, 356.3622, 347.48447, 338.84415, 330.3224, 321.8399, 313.43634, 305.03244, 296.7075, 288.69937, 280.61163, 272.52356, 264.4352, 256.1879, 248.01959, 240.00957, 232.31647, 224.46446, 216.8501, 208.83887, 200.82732, 192.9741, 184.96193, 177.02878, 169.13498, 161.43924, 153.7432, 146.36426, 139.2231, 132.24037, 125.01937, 117.95682, 111.21145, 104.62459, 98.59306, 92.40262, 85.97389, 79.78307, 73.75081, 67.639, 61.60638, 55.652966, 49.461227, 43.50746, 37.751987, 32.43299, 27.272638, 22.350334, 17.189728, 11.7908, 5.9947343, 2.1835327, NaN, NaN, 501.2844, 496.61105, 490.4326, 482.19434, 474.03497, 465.8753, 457.63608, 449.3173, 441.07742, 432.99567, 424.83438, 416.67273, 408.66928, 400.824, 393.05768, 385.29108, 377.44492, 369.4399, 361.35538, 353.34976, 345.22495, 337.06018, 329.05362, 321.28458, 313.59454, 305.9042, 298.2136, 290.20554, 282.27646, 274.26776, 266.1002, 257.61505, 249.12958, 240.80237, 232.31621, 224.22626, 216.21532, 208.3627, 200.27182, 192.33926, 184.44608, 176.67157, 169.21413, 162.07376, 155.0125, 147.6336, 140.3338, 133.19243, 126.28887, 119.54379, 112.95721, 106.291046, 100.021484, 93.354904, 87.084946, 81.68787, 76.37002, 70.65516, 64.70202, 58.51056, 53.073036, 47.91321, 42.83264, 38.30765, 33.22684, 27.828342, 22.747272, 18.06305, 13.219927, 7.0269146, 3.056936, NaN, NaN, 501.16492, 496.88763, 491.02603, 483.50076, 476.21286, 468.60782, 461.08173, 453.55536, 445.87027, 438.10565, 430.2615, 422.41705, 414.17612, 406.01407, 398.08945, 389.84753, 381.68454, 373.3627, 365.35757, 357.4314, 349.30676, 340.9836, 332.26376, 323.62283, 314.98154, 306.02274, 297.46, 289.37262, 280.88846, 272.95905, 265.5051, 258.1302, 250.755, 243.22095, 235.68661, 228.38994, 220.93439, 213.39923, 205.62585, 198.01082, 190.43517, 183.05756, 175.67967, 168.30154, 160.76447, 153.30644, 145.61012, 137.99286, 130.29597, 123.15426, 116.48844, 110.13984, 103.711685, 97.045235, 90.7754, 84.58474, 78.79075, 72.837845, 66.646645, 60.61401, 54.81934, 49.10389, 43.467663, 37.990055, 32.750465, 26.796225, 21.079992, 16.078156, 10.838007, 5.597724, 2.104127, NaN, NaN, 501.12473, 496.60983, 490.74823, 482.4308, 474.19226, 465.71573, 457.00116, 448.68237, 440.44247, 431.6476, 422.9316, 414.53223, 405.89474, 397.33615, 389.01495, 380.45566, 371.81677, 363.336, 354.30008, 345.73935, 337.1386, 328.4979, 319.93607, 311.29465, 302.8114, 294.4864, 286.3989, 278.4697, 270.77808, 262.76895, 254.91815, 246.90842, 238.89838, 230.88803, 222.5601, 214.15251, 205.66527, 197.09834, 188.68973, 180.04276, 172.06978, 163.89815, 156.1229, 148.50603, 141.36496, 134.1443, 126.92338, 119.543495, 112.32207, 105.6559, 98.91016, 92.00546, 85.73548, 79.78278, 73.909294, 67.71813, 61.84429, 56.52594, 51.20745, 46.206356, 40.609753, 35.052685, 29.65425, 24.33506, 19.174522, 13.934459, 7.90028, 3.3745286, NaN, NaN, 500.09454, 495.73804, 489.8764, 482.11346, 474.271, 466.2698, 458.26828, 450.42493, 442.34357, 434.18268, 426.3384, 418.41458, 410.1735, 402.1698, 394.24506, 386.39926, 378.39465, 370.78604, 363.49417, 356.12277, 348.4737, 340.70544, 333.01614, 325.32657, 317.71597, 310.02582, 302.17682, 294.48608, 286.95364, 279.18307, 271.3329, 263.5617, 255.6316, 247.70123, 239.84984, 231.76022, 223.90823, 216.05594, 208.12402, 200.1918, 192.37827, 184.3661, 176.5123, 168.81686, 161.43849, 153.98051, 146.52228, 138.90506, 131.52562, 124.30462, 117.08336, 110.338, 103.671776, 96.76725, 90.65615, 84.782974, 78.90963, 72.55988, 66.44806, 60.812325, 55.45426, 49.818222, 44.578945, 39.815853, 34.7351, 29.892387, 24.890778, 19.571472, 14.093237, 8.297262, 3.2951255, NaN, NaN, 501.28204, 496.68796, 490.50952, 481.6376, 472.44843, 463.25882, 454.14804, 445.3538, 436.6384, 427.9226, 419.12726, 410.5692, 402.32782, 394.0861, 385.84406, 377.5224, 369.51746, 361.3537, 353.50665, 345.58005, 337.85132, 329.9241, 322.07587, 314.06876, 306.2199, 298.21222, 290.28348, 282.03726, 274.0286, 265.78174, 257.85178, 249.84216, 241.75294, 233.5841, 225.41493, 217.40407, 209.55154, 201.6987, 193.9249, 186.1508, 178.57474, 171.03806, 163.65977, 156.36057, 149.37848, 142.39615, 135.25488, 127.87532, 120.73355, 113.75025, 107.32223, 100.973366, 94.465576, 87.95758, 81.76686, 75.73469, 69.464226, 63.27294, 57.24023, 51.604244, 46.444405, 40.72874, 35.092304, 29.45571, 23.977745, 18.896603, 13.815335, 8.416349, 3.493621, NaN, NaN, 502.66742, 498.4694, 493.0039, 485.87482, 478.9039, 471.299, 463.2977, 455.13766, 446.58115, 438.26196, 429.784, 421.2264, 412.90622, 404.18945, 395.9478, 387.4681, 379.3843, 371.3002, 363.295, 355.28955, 347.363, 339.19836, 331.11267, 323.18524, 315.0989, 307.25012, 299.32175, 291.31378, 283.2262, 274.90042, 267.1294, 259.59598, 252.06229, 244.3697, 236.67683, 228.98367, 221.36954, 213.59648, 205.82315, 197.81154, 189.7996, 181.8667, 174.01282, 166.3173, 158.85954, 151.16347, 143.54645, 136.24654, 129.34312, 122.36012, 115.059456, 107.8379, 100.7748, 94.26702, 87.91776, 81.568306, 75.21866, 68.78944, 62.201256, 55.851006, 49.937157, 44.142212, 38.66465, 33.34572, 28.185425, 23.342573, 18.42021, 13.49773, 8.1781435, 3.4936156, NaN, NaN, 501.51813, 496.76562, 490.42877, 482.03217, 473.87286, 465.5548, 457.07797, 448.60077, 439.88553, 431.40762, 422.85013, 414.2923, 405.49637, 396.7793, 387.90338, 379.10632, 370.38815, 361.66962, 353.34702, 344.7863, 336.42337, 328.09976, 319.37946, 310.4209, 301.3827, 292.42334, 283.7015, 274.9, 266.4153, 258.00955, 249.92068, 242.38666, 234.69373, 226.92119, 219.14836, 211.61319, 204.15707, 196.54202, 188.76805, 181.39043, 174.09189, 166.79308, 159.33533, 151.8773, 144.65704, 137.27785, 130.13643, 123.391525, 116.487686, 109.66298, 102.67932, 95.85415, 89.26685, 82.599976, 75.77414, 69.186195, 62.836174, 56.803467, 50.53244, 44.89629, 39.259983, 34.020462, 28.939585, 24.096758, 19.333208, 14.648944, 9.805778, 4.8830976, 1.548312, NaN, NaN, 499.8542, 495.02246, 488.68558, 479.8136, 471.17892, 461.9893, 452.95773, 443.60886, 434.73495, 425.7022, 416.43134, 407.16003, 398.20532, 389.48798, 380.69098, 372.05215, 363.72998, 355.32822, 346.92612, 339.07855, 330.9929, 322.8276, 314.8206, 306.5754, 298.25058, 290.1633, 281.99643, 273.9085, 265.82028, 257.89032, 249.80145, 241.87088, 233.78139, 225.53294, 217.83939, 209.82828, 202.13412, 194.59834, 186.90363, 179.1293, 171.35466, 163.57974, 155.88387, 148.42574, 141.12602, 133.82603, 126.44646, 119.22531, 111.8452, 104.782265, 97.87781, 91.36995, 84.861885, 78.353615, 71.52764, 64.86019, 58.58942, 52.556595, 46.99989, 41.125492, 35.409702, 30.011309, 24.850948, 19.928637, 14.76802, 9.527877, 4.2082005, 1.3498095, NaN, NaN, 499.97232, 495.69504, 489.83347, 482.14978, 474.94113, 467.33612, 459.88925, 452.20447, 444.36093, 436.43787, 428.51447, 420.51157, 412.74606, 404.90103, 397.21417, 389.52704, 381.99814, 374.31042, 366.54318, 358.85492, 351.16635, 343.87384, 336.73962, 329.68442, 322.47043, 315.2562, 307.88312, 300.5098, 292.81906, 285.04874, 277.19882, 269.50723, 261.9739, 254.44034, 246.9858, 239.53098, 231.91727, 224.30327, 216.76831, 209.31241, 201.73723, 194.20145, 186.82404, 179.36703, 171.9891, 164.53156, 157.07375, 149.77435, 142.55405, 135.65086, 129.14423, 122.3993, 115.73352, 109.226234, 102.56002, 95.6555, 88.909485, 82.163246, 75.49615, 69.22571, 63.153522, 57.51773, 51.723026, 45.928158, 40.37128, 34.89364, 29.098291, 23.382174, 18.062864, 12.6640215, 7.265036, 2.8187058, NaN, NaN, 498.9418, 494.18927, 488.2484, 480.32706, 472.72226, 465.03793, 457.27414, 449.4308, 441.4287, 433.58478, 425.50284, 417.49982, 409.65497, 401.57208, 393.40964, 385.3261, 377.4008, 369.31665, 361.15292, 353.1474, 345.02267, 336.62018, 328.13806, 319.57632, 310.93494, 302.45175, 293.80966, 285.2465, 276.84155, 268.43628, 260.18924, 252.0212, 244.01143, 235.76343, 227.83234, 219.82164, 211.81061, 203.64064, 195.70831, 187.77568, 180.08073, 172.46483, 164.84865, 157.31151, 149.85345, 142.55382, 135.17456, 127.71569, 120.41526, 113.74943, 107.24209, 100.81391, 94.06807, 87.401375, 80.97257, 74.94043, 69.2256, 63.034355, 56.9223, 51.206966, 45.570858, 40.410904, 35.488983, 30.56694, 25.247828, 20.484325, 15.641316, 10.560005, 5.5579653, 2.1438046, NaN, NaN, 499.0597, 494.22797, 487.9703, 479.49442, 470.93896, 462.1455, 453.27246, 444.39902, 436.00058, 427.52255, 419.20267, 410.80322, 402.56192, 394.08252, 385.9198, 377.836, 369.83115, 361.826, 353.74124, 345.6562, 337.33298, 329.00946, 320.52704, 312.04428, 303.5612, 295.157, 286.91107, 278.74408, 270.73538, 262.40915, 254.32051, 246.39015, 238.22157, 229.97334, 221.80411, 213.95181, 206.17854, 198.24632, 190.47246, 182.69829, 175.2015, 167.58543, 159.88974, 152.4318, 145.29094, 138.22919, 130.92915, 123.7082, 116.56635, 109.58297, 102.59935, 95.61549, 89.02823, 82.28201, 75.77369, 69.82077, 63.867683, 58.073177, 52.51665, 47.515644, 42.31606, 37.55296, 32.472202, 26.200466, 20.56368, 14.212185, 7.3841076, 2.4613988, NaN, NaN, 498.6628, 493.59344, 487.25656, 479.09753, 471.25504, 462.93695, 454.6185, 446.5374, 438.37677, 430.29504, 422.3715, 414.36838, 406.44418, 398.8367, 390.9119, 383.14532, 375.1407, 367.215, 359.44754, 351.91757, 343.9117, 336.0641, 327.97836, 320.13013, 312.36087, 304.59134, 296.66293, 289.0514, 281.43954, 273.66882, 265.65994, 257.80933, 250.19633, 242.50375, 235.04881, 227.5143, 219.58292, 211.65123, 203.87788, 196.02492, 188.64761, 181.27005, 173.81288, 166.43478, 159.69113, 152.55054, 145.72708, 138.98274, 132.0795, 125.176, 118.5897, 111.84447, 105.178375, 98.59143, 92.32173, 86.21057, 80.41671, 74.62268, 68.987236, 63.748512, 58.350903, 52.71501, 47.158344, 41.522144, 36.679653, 32.233982, 27.70883, 22.38966, 16.99096, 12.544863, 7.1459026, 2.6201932, NaN, NaN, 498.66205, 493.67188, 487.49344, 478.6215, 469.43228, 460.24268, 451.36957, 442.33762, 433.54294, 424.82715, 416.19025, 407.55295, 398.83606, 390.67355, 382.66922, 374.66458, 366.81815, 358.7336, 350.72806, 342.4051, 334.2007, 325.95636, 317.71167, 309.3081, 301.30063, 293.29282, 285.2847, 277.59344, 269.7433, 262.13077, 254.43863, 246.66692, 238.49837, 230.40881, 222.23961, 213.99077, 205.74161, 198.04736, 190.67015, 183.29266, 176.15292, 169.01292, 161.63466, 154.01811, 146.71866, 139.33958, 132.1983, 124.89808, 117.83565, 110.93169, 104.10686, 97.51988, 91.01207, 84.424675, 77.757706, 71.01114, 64.581856, 58.46988, 52.67524, 47.11858, 41.442696, 35.96512, 30.566786, 25.088919, 19.610905, 14.7679, 10.321763, 5.00215, 1.9055954, NaN, NaN, 499.77014, 495.09686, 488.83926, 481.0764, 473.6301, 465.70822, 457.54837, 449.1505, 441.06924, 433.06686, 424.90573, 416.98196, 409.05792, 401.45053, 393.92212, 386.4727, 378.78522, 371.01822, 363.25092, 355.3248, 347.2002, 338.71857, 330.39514, 322.3885, 314.4608, 306.69135, 298.68378, 290.67587, 282.58838, 274.57986, 266.17453, 258.16537, 250.2352, 242.38403, 234.53256, 226.83942, 219.38394, 212.00749, 204.6308, 197.33315, 189.51962, 181.66612, 174.12967, 166.5136, 158.5799, 150.16982, 142.15614, 134.45953, 127.08004, 119.70028, 112.55833, 105.09869, 98.03558, 91.2897, 84.464226, 77.956, 71.3682, 65.17706, 58.826984, 52.714844, 47.118507, 41.085403, 35.131508, 29.65377, 24.49345, 19.174215, 14.01363, 8.535328, 3.7714677, NaN, NaN, 499.45248, 494.93762, 488.91763, 480.6795, 472.67868, 464.28146, 455.88388, 447.3275, 438.6916, 430.1345, 421.73553, 413.41547, 404.93658, 396.3781, 387.97778, 379.49786, 370.93832, 362.29916, 353.81818, 345.1783, 336.61734, 327.8182, 319.33582, 311.09088, 302.6078, 294.20364, 286.1163, 278.2665, 270.25784, 262.24884, 254.08095, 245.99202, 237.66486, 229.7339, 221.64403, 213.39519, 205.14603, 197.21382, 189.36064, 181.42783, 173.61371, 165.91829, 158.2226, 150.60594, 142.90967, 135.45114, 128.30975, 120.77135, 112.99459, 105.05883, 97.67829, 91.1705, 84.34503, 77.836815, 71.16965, 64.264145, 57.199646, 50.92871, 45.054493, 39.497646, 33.900955, 28.264418, 22.627726, 17.149664, 11.274478, 4.0493555, NaN, NaN, 500.71875, 496.36237, 490.7385, 483.68863, 476.797, 469.19214, 461.50778, 453.98157, 446.1382, 438.61145, 430.92596, 423.63635, 416.26724, 408.81866, 401.5283, 393.92065, 386.2335, 378.54605, 370.46204, 362.13992, 353.7382, 345.09836, 336.7752, 328.13464, 319.81082, 311.48666, 303.16217, 294.9959, 286.98788, 279.13815, 271.44672, 263.83426, 256.22156, 248.37064, 240.51942, 232.74722, 224.7368, 217.04332, 209.27022, 201.7348, 193.92148, 186.30617, 178.7699, 171.3127, 164.09323, 157.19087, 150.20892, 143.22676, 136.165, 129.10298, 122.19945, 115.53374, 108.94717, 102.51911, 96.09084, 89.662384, 83.07498, 76.408, 70.05829, 64.34338, 58.62832, 52.992474, 46.959568, 40.847095, 35.369534, 30.0506, 24.9697, 20.365025, 15.522063, 10.520197, 5.359413, 1.6276885, NaN, NaN, 499.6882, 494.85654, 488.67816, 480.2024, 471.3302, 462.4576, 453.18854, 443.60214, 434.3322, 425.22034, 415.87033, 406.59915, 397.64456, 389.00656, 380.6852, 372.36353, 364.2, 356.0362, 347.9513, 339.46976, 331.10678, 322.7038, 313.9041, 305.10403, 296.38287, 287.81992, 279.3359, 270.93082, 262.4461, 254.04033, 245.71352, 237.30707, 228.90027, 220.49313, 212.32361, 203.9951, 195.90424, 187.73373, 179.5629, 171.39174, 163.45825, 155.52448, 147.74907, 140.3701, 132.99086, 125.61135, 118.23158, 111.01026, 103.471245, 96.328766, 89.503494, 83.07484, 76.64597, 70.45503, 64.34328, 58.390087, 52.43673, 46.562576, 40.92641, 35.845787, 30.68565, 25.604774, 20.44438, 15.045674, 9.885014, 4.7242227, 1.8658825, NaN, NaN, 499.0144, 493.70746, 487.6875, 479.29092, 470.9732, 462.4175, 454.01993, 445.4635, 437.06522, 428.82504, 420.4261, 411.78903, 402.5177, 393.48367, 384.84552, 376.0485, 367.33032, 359.00812, 350.68555, 342.36267, 334.03946, 325.55734, 317.23343, 308.67136, 300.50534, 292.339, 284.25162, 276.08463, 267.9173, 259.82898, 251.81961, 243.65134, 235.72066, 227.39311, 219.14455, 211.1336, 203.36032, 195.50742, 187.49554, 179.5627, 171.43121, 163.41841, 155.48463, 148.02661, 140.56831, 132.95103, 125.57154, 118.19178, 110.73239, 103.59017, 96.76515, 90.01927, 83.035065, 76.60621, 70.3359, 64.224144, 58.19158, 52.317604, 46.28469, 40.17222, 34.29772, 28.89939, 24.294815, 19.293177, 13.815052, 7.9397993, 3.1759567, NaN, NaN, 499.29105, 494.38016, 488.2018, 479.80527, 471.40836, 462.93192, 454.4551, 445.81952, 437.342, 428.86417, 420.386, 412.14514, 404.14172, 396.21725, 388.3717, 380.7636, 373.5515, 366.33917, 358.8888, 351.43817, 344.0665, 336.9324, 329.32242, 321.71216, 314.10162, 306.49078, 298.6418, 291.1097, 283.57733, 276.20325, 268.51172, 261.0578, 253.6036, 246.38705, 239.24957, 231.79459, 224.41866, 216.72519, 208.8728, 201.17876, 193.64307, 186.02779, 178.33287, 170.47902, 163.02155, 155.24644, 147.47104, 139.69534, 132.07806, 124.14308, 116.04908, 108.351555, 101.36798, 94.62226, 88.03504, 81.44762, 75.09809, 68.98649, 63.192196, 57.397747, 51.761887, 45.967113, 40.172173, 34.456455, 29.216908, 23.897837, 18.816803, 13.815036, 8.57496, 3.5729437, NaN, NaN, 500.51794, 495.84473, 489.5872, 480.87384, 472.16016, 463.28766, 454.494, 445.8584, 437.14322, 428.66537, 420.26642, 411.7879, 403.38824, 395.0675, 386.82568, 378.42505, 370.1033, 362.17752, 354.2514, 346.1665, 337.8038, 329.5597, 321.236, 312.83264, 304.3497, 295.7078, 287.22415, 278.81943, 270.57294, 262.32614, 253.9204, 245.51431, 237.42511, 229.4149, 221.56302, 213.71083, 205.85834, 198.00554, 190.23178, 182.53705, 174.80235, 166.94838, 158.93542, 151.3982, 143.78136, 136.32292, 129.10226, 121.881355, 114.342766, 106.96262, 99.82029, 92.51898, 85.29678, 78.39181, 71.96282, 65.69238, 59.024876, 52.198387, 45.927345, 39.735497, 33.980083, 28.184814, 22.865723, 17.864065, 13.259255, 8.733738, 4.0493245, NaN, NaN, 501.30914, 496.79437, 490.69528, 482.9326, 475.2488, 467.08942, 458.9297, 450.9281, 442.847, 434.76556, 426.60458, 418.44327, 409.88544, 401.56497, 393.32343, 385.1608, 377.0771, 369.38934, 361.46356, 353.37894, 345.65067, 337.8825, 329.9555, 321.7111, 313.54562, 305.5384, 297.45157, 289.44373, 281.59412, 273.74423, 265.97336, 258.12286, 250.11348, 242.3417, 234.64894, 226.95589, 219.10391, 211.25163, 203.31975, 195.46687, 187.85167, 180.47418, 173.17577, 165.55974, 158.02277, 150.2475, 142.47194, 134.69609, 127.07863, 119.4609, 111.4461, 103.58971, 96.28855, 88.8284, 81.76482, 75.01847, 68.35127, 61.04886, 54.38121, 47.951485, 41.95816, 35.7662, 29.812218, 23.93745, 18.459475, 13.219536, 7.9000654, 3.0568454, NaN, NaN, 499.05112, 494.3779, 488.19955, 479.80304, 471.24774, 462.61288, 453.9777, 445.26288, 436.62692, 427.75293, 418.72006, 410.3207, 401.8418, 393.44177, 385.19992, 376.87848, 368.7152, 360.5516, 351.99136, 343.74786, 335.58328, 327.5769, 319.6495, 311.64255, 303.47668, 295.78622, 288.01617, 280.16653, 272.3959, 264.70425, 257.09164, 249.71666, 242.10347, 234.80725, 227.59007, 220.53128, 213.47224, 206.49228, 199.35342, 192.21434, 184.99567, 177.69742, 170.24023, 162.94145, 155.64241, 148.58115, 141.36095, 134.21983, 126.91977, 119.61945, 112.31887, 104.7006, 96.764595, 89.383835, 82.24091, 75.256485, 68.27181, 61.763157, 55.492428, 48.983364, 42.712242, 36.5997, 30.963295, 25.564905, 19.769415, 14.132547, 8.892503, 4.0493126, 1.4291784, NaN, NaN, 499.80307, 495.12985, 489.10995, 481.42642, 474.2971, 466.69223, 459.08707, 451.24396, 443.4798, 435.7153, 427.6336, 419.15543, 410.83536, 402.4357, 394.0357, 385.3184, 376.60068, 367.96188, 359.5605, 351.238, 343.0341, 335.02805, 327.02167, 318.8564, 311.008, 303.00067, 295.1516, 287.38156, 279.6112, 271.76126, 263.67313, 255.66399, 247.57521, 239.64474, 231.63466, 223.8622, 215.85149, 207.9198, 199.82915, 191.97617, 184.47984, 177.02292, 170.12105, 163.37762, 156.23729, 149.33473, 142.3526, 135.21152, 128.2289, 121.3254, 114.65972, 107.993835, 101.089645, 94.264595, 87.59804, 80.93127, 74.66113, 68.232056, 62.040905, 56.246452, 50.689976, 45.530254, 40.05287, 34.17841, 28.303782, 22.825935, 17.427336, 11.869804, 7.503067, 3.2950315, NaN, NaN, 498.69348, 494.09943, 488.15872, 480.0791, 472.07837, 463.76044, 455.36298, 447.1236, 439.04236, 430.88156, 422.95816, 415.03445, 407.26892, 399.42386, 391.65775, 383.97058, 376.3624, 368.67465, 360.74887, 352.82278, 344.65857, 336.17697, 327.93283, 320.00546, 312.15707, 304.14984, 296.22156, 288.37225, 280.52264, 272.67276, 264.66397, 256.57556, 248.32825, 240.08058, 231.7533, 223.42566, 215.177, 207.08665, 199.23396, 191.38095, 183.68631, 175.99138, 168.37549, 160.75931, 153.14285, 145.28809, 137.51236, 129.9744, 122.43615, 115.056335, 107.75561, 100.772064, 93.788284, 87.04236, 80.53432, 73.94669, 67.43823, 60.92957, 54.341316, 48.149754, 42.394608, 36.996532, 31.518927, 26.120564, 20.642666, 15.323409, 9.686434, 5.160862, 2.2231565, NaN, NaN, 487.20752, 481.90033, 475.48398, 466.2948, 457.026, 448.07367, 439.2002, 430.4848, 421.9275, 413.29062, 404.41565, 395.778, 387.21927, 378.6602, 370.33853, 362.0165, 353.3771, 344.97513, 336.81064, 328.48727, 319.92575, 311.5224, 303.19803, 295.2697, 287.2618, 279.09503, 270.92792, 262.44327, 253.879, 245.47298, 237.46313, 229.6116, 222.07703, 214.30423, 206.45181, 198.67842, 190.98405, 183.28941, 175.4358, 167.8199, 160.2434, 152.54759, 145.01018, 137.4725, 130.01389, 122.71371, 115.41326, 108.27128, 101.12904, 94.22464, 87.399376, 80.494514, 73.74816, 67.00159, 60.334167, 53.269638, 46.125484, 39.536766, 33.265377, 26.914412, 20.682333, 13.854615, 7.42365, 2.977432, NaN, NaN, 382.22614, 377.31253, 371.05145, 362.17465, 353.13898, 344.18216, 335.14566, 326.6637, 318.4192, 310.0158, 301.6121, 293.04944, 284.2486, 275.76453, 267.2801, 258.79532, 250.1516, 241.5075, 233.10098, 224.45618, 215.85066, 207.52242, 199.03517, 190.78555, 182.53561, 174.28534, 166.27274, 158.25981, 150.16724, 141.91566, 133.98114, 126.284355, 118.98405, 112.0009, 105.09688, 98.51006, 91.76431, 85.0977, 78.668976, 71.92257, 65.21563, 58.548157, 52.436115, 46.40327, 40.211483, 34.098896, 27.74796, 21.238047, 15.204284, 8.37639, 2.7392364, NaN, NaN, 321.19363, 316.5164, 310.25348, 302.00833, 293.76285, 285.51703, 277.42947, 269.73807, 262.12567, 254.43372, 246.58284, 238.33514, 229.53194, 221.04562, 212.79689, 204.30988, 195.26724, 186.1449, 177.57745, 169.40631, 161.11584, 152.86472, 144.45456, 136.20276, 128.10931, 120.015564, 111.842125, 103.66837, 95.17684, 87.47861, 80.01819, 72.954346, 66.04901, 59.14344, 51.999504, 44.617172, 37.47273, 30.010485, 23.18309, 16.990604, 10.480352, 4.0492907, NaN, NaN, 264.7424, 261.01547, 255.86105, 247.85164, 239.76259, 231.356, 223.50426, 216.04878, 208.51372, 200.2645, 192.25291, 184.47899, 176.54613, 168.85094, 160.83813, 152.82501, 144.73222, 136.08371, 127.990265, 119.7378, 112.00082, 104.1445, 96.60532, 88.74842, 80.89121, 72.95433, 64.8584, 56.524014, 48.26867, 41.04497, 33.741634, 26.358644, 19.451738, 13.100353, 5.3196387, 1.5879663, NaN, NaN, 208.98962, 204.58743, 198.87636, 190.42844, 181.86118, 173.41254, 165.32057, 156.75226, 147.58853, 137.71028, 127.47449, 116.76206, 105.69197, 94.621284, 84.50239, 75.21637, 66.40617, 58.66717, 51.40415, 44.379017, 37.869637, 31.439438, 25.723536, 20.325037, 14.3706455, 8.019103, 2.7789328, NaN, NaN, 197.32957, 192.72884, 186.54147, 177.49806, 168.2956, 159.41006, 150.28612, 141.00308, 131.95767, 122.59445, 113.0721, 103.311226, 93.47053, 83.867455, 74.97826, 66.48554, 57.913094, 49.975327, 42.196014, 34.733948, 27.192219, 20.285341, 13.775196, 7.34424, 2.1834502, NaN, NaN, 190.98369, 186.46213, 180.3539, 172.02422, 163.45618, 154.72911, 146.08102, 137.35321, 128.46634, 119.49972, 110.532715, 101.8034, 92.676895, 83.15315, 73.708336, 64.501205, 55.690544, 47.35579, 39.33823, 31.955444, 24.493004, 17.268469, 9.964283, 3.136221, NaN, NaN, 195.46545, 190.70602, 184.75658, 177.2997, 169.92189, 161.75044, 153.26132, 144.53383, 135.72661, 127.15706, 118.58715, 110.01689, 101.60499, 93.748276, 85.8119, 78.58952, 71.84312, 65.33462, 58.90528, 52.078854, 44.73622, 37.11548, 29.256292, 21.634974, 13.140046, 4.4859715, NaN, NaN, 191.61824, 186.70007, 180.11588, 171.07219, 162.10744, 153.1423, 144.33545, 135.68692, 126.879326, 118.07135, 109.10429, 99.9781, 91.168976, 82.35947, 73.70832, 65.13618, 56.643055, 47.75268, 38.623768, 29.097515, 20.32503, 12.703381, 4.366876, NaN, NaN, 188.4452, 183.28899, 176.38736, 167.26418, 158.21992, 149.09595, 139.8922, 130.37065, 120.84866, 111.16753, 101.80336, 93.07367, 84.50234, 76.3275, 68.39045, 60.77059, 53.229824, 46.40321, 39.496983, 32.193592, 24.215134, 16.196669, 7.8603086, 2.1437504, NaN, NaN, 192.60974, 187.53294, 181.50409, 173.17444, 164.84447, 156.67284, 148.65955, 140.16989, 131.91792, 123.66562, 115.33363, 106.52516, 98.271835, 90.09755, 82.63723, 75.25601, 68.19201, 61.365894, 54.53955, 47.79236, 41.12433, 34.05915, 26.993734, 20.642588, 13.735492, 5.3990316, 1.111577, NaN, NaN, 193.6806, 189.87303, 184.79617, 177.41862, 169.96149, 162.02806, 154.253, 146.39832, 138.38463, 130.37064, 122.27697, 114.500404, 106.80291, 99.26384, 92.04194, 84.81979, 77.51802, 69.8985, 62.278698, 54.420483, 46.998554, 39.695435, 32.07451, 24.21513, 17.149372, 9.289421, 2.778931, NaN, NaN, 186.85866, 181.74205, 174.8404, 165.32047, 155.80011, 146.04128, 135.32982, 124.73684, 114.14331, 103.78731, 93.311745, 83.549934, 75.09727, 66.763306, 58.54807, 50.3325, 41.759384, 33.42407, 25.326576, 16.990587, 8.49547, 2.461341, NaN, NaN, 183.05096, 177.65662, 170.91347, 161.79005, 152.82489, 144.3354, 136.16295, 128.38692, 120.68994, 113.230736, 106.48547, 99.89871, 93.153015, 85.77218, 78.3117, 70.692215, 63.310562, 56.722412, 50.53095, 45.053726, 39.536667, 33.582836, 27.390673, 20.642586, 13.497311, 6.1929946, 1.5879651, NaN, NaN, 186.8983, 181.54372, 174.88004, 166.07413, 156.91083, 147.27106, 137.27379, 127.276024, 116.80165, 106.20772, 95.73228, 85.73249, 76.44653, 67.39828, 58.82588, 50.491253, 42.39444, 34.773613, 27.390669, 20.24563, 12.822466, 4.8035564, NaN, NaN, 184.59781, 179.28284, 171.50844, 162.70238, 154.13396, 145.40651, 136.99606, 128.50592, 120.174126, 111.92136, 103.74761, 95.097374, 86.52613, 77.79579, 69.06509, 60.651505, 51.76131, 42.63258, 33.820988, 25.644125, 18.260853, 9.44821, 2.6201355, NaN, NaN, 176.66493, 171.9844, 165.79642, 157.54549, 149.13554, 140.56656, 132.07657, 123.58622, 115.09553, 106.68384, 98.11308, 89.78006, 81.208595, 72.3193, 63.429607, 54.777664, 45.72845, 36.440685, 27.470053, 18.975372, 10.639129, 3.7316976, NaN, NaN, 166.15341, 160.67928, 153.53888, 144.33534, 135.76616, 127.11728, 118.468025, 109.73905, 101.32714, 92.756165, 84.10546, 75.53376, 66.64422, 58.230537, 50.21341, 42.19597, 34.73391, 27.747906, 21.238005, 14.966076, 7.701513, 2.223147, NaN, NaN, 165.20137, 160.20323, 153.45952, 143.85927, 134.25858, 124.73677, 115.6113, 106.644135, 97.755936, 88.708626, 79.66091, 70.850914, 62.199287, 53.388542, 44.33927, 35.448368, 26.398306, 18.22115, 10.4406395, 5.041744, 3.8507922, 3.9301891, NaN, NaN, 160.52055, 155.16528, 148.0247, 138.02747, 128.50584, 119.102806, 110.29451, 101.48583, 93.27199, 85.29592, 77.200485, 69.22379, 61.246784, 53.269463, 45.291836, 37.552048, 30.169209, 22.309765, 15.045464, 7.7809057, 2.461339, NaN, NaN, 155.40329, 150.16689, 143.10548, 133.98082, 124.69707, 115.17483, 106.04893, 97.55751, 89.1451, 80.97046, 72.63674, 64.22331, 55.809536, 47.474796, 39.298485, 31.439392, 23.579996, 16.037868, 8.892439, 5.081441, 4.088982, NaN, NaN, 158.06108, 153.5388, 147.42961, 138.46384, 129.49768, 120.68983, 111.08804, 101.56517, 92.51803, 83.31176, 73.946335, 64.89798, 56.2461, 47.4351, 39.179405, 31.47908, 23.540298, 16.156956, 9.4879, 3.295011, NaN, NaN, 158.10074, 153.41978, 147.3106, 138.90024, 130.9656, 123.189384, 115.09545, 106.92184, 98.98598, 91.20854, 83.58954, 76.367096, 68.50943, 60.25458, 51.602512, 42.71193, 33.582806, 24.453274, 16.037867, 8.813043, 5.637215, 5.1608367, NaN, NaN, 149.1751, 144.09723, 137.43234, 128.62483, 119.65823, 110.77061, 102.04131, 93.23228, 85.21653, 77.041725, 69.18408, 61.72301, 54.579178, 46.720673, 38.385567, 30.288279, 22.270061, 14.569102, 6.0738935, 1.1512748, NaN, NaN, 153.7768, 148.85773, 142.66905, 134.97261, 127.275894, 118.388596, 109.421555, 100.6922, 91.96248, 83.54984, 75.37498, 67.04103, 58.706753, 50.76903, 42.51347, 33.781265, 25.286854, 16.87148, 8.932134, 4.9623446, 3.930187, NaN, NaN, 147.6676, 142.11363, 135.60738, 127.27588, 119.26146, 111.08801, 102.67617, 94.58142, 86.56573, 79.02592, 71.80332, 64.34235, 56.246086, 47.43509, 38.22679, 29.018084, 19.967741, 10.996393, 2.8980236, NaN, NaN, 148.38168, 143.54182, 137.35298, 128.70418, 119.97564, 111.64352, 103.23169, 94.89888, 86.248276, 77.27983, 68.23162, 59.34176, 50.53089, 41.79903, 33.066795, 24.492966, 15.204244, 5.915101, 2.3422418, NaN, NaN, 142.43102, 137.1943, 130.76723, 122.27683, 113.23061, 104.66013, 96.0893, 87.51811, 78.78783, 69.9778, 61.72301, 53.944157, 46.40315, 39.020634, 31.796621, 24.572353, 17.427225, 9.090924, 2.4216394, NaN, NaN, 144.89067, 140.13007, 133.78244, 124.89542, 115.76996, 106.72344, 97.7559, 89.18477, 80.53392, 72.20019, 63.548622, 54.97607, 46.561916, 38.306187, 30.447056, 22.349455, 14.410318, 6.94725, 3.1362164, 2.1040492, NaN, NaN, 140.96318, 136.2025, 130.25148, 122.47523, 115.01609, 106.92184, 98.747894, 90.73236, 83.03397, 74.93845, 67.1601, 59.381454, 51.602512, 43.743893, 35.805584, 27.708197, 19.689878, 11.909427, 4.6050606, NaN, NaN, 139.41597, 134.53624, 127.99005, 118.34894, 108.11219, 97.39877, 87.39908, 77.87511, 68.82692, 59.77833, 50.729347, 41.799038, 32.63018, 23.579994, 14.648498, 7.026646, 3.2156136, 1.905555, NaN, NaN, 136.2025, 131.52104, 125.01444, 115.57157, 105.8902, 96.684525, 87.71654, 79.22436, 70.8112, 62.55645, 54.14261, 45.56966, 36.996353, 29.295946, 21.9922, 14.291229, 6.2723846, 2.7789283, NaN, NaN, 136.67857, 132.63191, 127.39493, 120.13435, 112.63546, 103.82689, 94.06559, 83.946686, 73.70822, 63.58831, 53.586964, 45.252136, 38.46495, 30.486748, 22.865486, 16.077562, 8.813043, 3.2156136, NaN, NaN, 134.37752, 129.25961, 122.8323, 113.429, 103.7872, 94.14494, 84.85938, 75.81151, 67.7157, 59.619576, 50.332447, 40.330456, 31.042452, 21.396772, 12.10791, 5.4387236, 2.5804343, NaN, NaN, 131.20361, 126.284004, 120.09465, 111.683174, 103.43007, 95.57344, 88.192696, 81.20852, 74.303474, 67.71569, 60.81019, 52.872547, 45.25212, 38.42525, 31.042446, 23.183039, 15.6409, 7.3045287, 3.0171194, NaN, NaN, 130.68784, 125.33179, 118.42823, 108.429565, 98.54945, 87.83554, 77.95443, 68.07285, 58.78611, 49.37988, 40.33044, 31.518757, 22.706697, 14.251526, 5.796005, 0.793983, NaN, NaN, 125.9269, 120.53105, 114.26217, 106.564674, 98.94624, 91.24818, 83.54981, 75.53368, 67.59661, 59.976738, 52.832848, 45.609325, 37.432945, 28.303589, 19.49139, 11.472754, 5.597514, 2.6598308, 2.1834457, NaN, NaN, 126.64104, 122.11807, 115.9286, 107.04081, 97.99391, 89.105354, 80.454506, 71.962036, 63.46921, 55.69043, 48.22887, 40.370125, 32.66985, 25.525007, 18.776869, 12.02851, 6.5502667, 4.1683755, 3.6919942, NaN, NaN, 126.76005, 121.68163, 114.85731, 105.969475, 97.0019, 87.79584, 78.82746, 70.09681, 60.968914, 52.158123, 43.029427, 34.059093, 25.882254, 18.57839, 10.718508, 3.8904865, NaN, NaN, 126.720345, 121.721275, 115.45243, 107.199486, 99.18429, 91.16877, 83.232315, 75.21617, 66.406, 57.357315, 48.30823, 39.655666, 31.24089, 23.22272, 16.077547, 9.408496, 5.359323, 3.374405, 3.2156105, NaN, NaN, 123.82403, 118.507484, 112.317894, 104.858406, 97.39864, 89.383064, 81.2878, 72.87474, 64.143845, 55.015686, 45.80774, 36.758152, 28.422647, 20.404367, 12.54456, 6.272376, 3.7316902, 3.0965135, NaN, NaN, 124.22073, 119.69772, 113.666885, 105.969376, 98.827095, 91.52584, 84.14496, 76.68445, 69.223656, 61.60385, 53.507496, 44.934536, 36.99629, 28.740187, 20.721922, 11.909407, 3.7316887, NaN, NaN, 122.23692, 117.55517, 111.2862, 102.398224, 92.95433, 83.66873, 75.17641, 66.604355, 57.714447, 48.50663, 39.457165, 30.88362, 22.627272, 14.529378, 6.9869337, 3.8110843, 3.0171142, NaN, NaN, 122.71299, 117.832855, 111.28616, 101.406204, 91.64481, 81.40676, 72.00159, 62.834106, 53.666214, 44.616978, 36.281807, 28.303535, 20.20587, 11.750611, 5.438711, 2.937716, 1.9849478, NaN, NaN, 117.23767, 112.23838, 106.445404, 98.43018, 90.3353, 82.16072, 74.144554, 66.048706, 57.3969, 48.903492, 40.72726, 33.027016, 25.485258, 17.943222, 10.003938, 3.0965092, NaN, NaN, 118.94371, 113.58737, 106.68344, 96.68423, 86.92262, 77.16055, 67.75519, 58.70658, 48.943165, 39.89373, 30.962973, 22.38908, 13.695739, 6.5502505, 3.8110805, 2.858317, NaN, NaN, 113.23024, 108.07214, 101.16803, 92.438354, 83.54957, 74.819145, 66.08835, 57.515926, 49.02253, 40.211246, 31.478973, 22.825714, 14.41027, 5.75629, 2.3422341, NaN, NaN, 109.421165, 104.104256, 97.358734, 87.59716, 77.67639, 67.75514, 58.46842, 49.101894, 39.655556, 30.923262, 22.42876, 14.25148, 5.2005157, NaN, NaN, 114.49984, 110.05598, 104.183586, 95.45404, 86.00984, 76.96206, 68.23135, 59.81778, 51.245102, 42.989594, 34.733753, 26.39819, 18.062286, 9.805439, 5.3593063, 3.3743944, 3.2949977, NaN, NaN, 109.897224, 105.05648, 98.94587, 90.37483, 82.041534, 74.26349, 67.19949, 60.294006, 53.22953, 45.76791, 38.385403, 30.605696, 22.508135, 14.727825, 7.502987, 4.4859457, 3.533187, NaN, NaN, 108.42911, 103.8264, 97.00151, 88.82722, 80.49386, 72.00143, 63.667385, 55.412384, 47.236427, 38.980762, 30.407219, 21.595148, 13.020877, 4.1286607, NaN, NaN, 107.15937, 101.6837, 94.70001, 85.57325, 76.366714, 67.239136, 57.9524, 48.824, 39.695194, 30.248438, 21.198193, 12.862087, 5.716583, 2.9377084, 1.9849427, NaN, NaN, 107.55612, 102.39789, 95.969765, 86.208145, 77.00164, 68.27095, 60.095512, 51.91975, 44.140564, 35.964165, 27.787436, 19.689774, 11.512396, 5.478393, 3.3346915, 2.7789135, NaN, NaN, 104.54052, 99.779015, 92.87463, 84.30336, 76.36667, 68.27093, 59.85737, 51.760975, 43.5055, 35.32908, 27.231716, 19.372206, 10.877243, 3.8904672, NaN, NaN, 105.492775, 100.57257, 94.223755, 86.049355, 77.7159, 69.77896, 61.52421, 53.42789, 44.85496, 36.281677, 27.70803, 19.134027, 10.877239, 5.08141, 2.9377055, 2.6995146, NaN, NaN, 102.715225, 97.318794, 90.255615, 81.20803, 71.92194, 63.270416, 54.777283, 45.966274, 36.5992, 27.072924, 18.181332, 8.971776, 3.5728784, 1.8261456, NaN, NaN, 105.175285, 100.017, 93.588806, 84.382645, 75.096695, 66.04845, 57.317303, 48.34765, 39.695133, 31.04225, 22.468391, 13.973565, 4.366842, NaN, NaN, 105.13557, 100.61216, 94.58079, 86.64451, 79.2635, 71.56473, 64.02442, 56.24571, 48.62546, 41.00493, 33.622265, 26.318724, 18.935532, 11.710861, 6.153248, 4.088953, 3.7713673, NaN, NaN, 99.85822, 95.17597, 89.14445, 80.73176, 72.00124, 63.111614, 54.221596, 45.489952, 36.916702, 28.581255, 20.245468, 12.147521, 6.4311304, 4.2080464, 3.6522717, NaN, NaN, 98.82652, 93.27128, 86.36669, 78.58883, 70.890045, 62.873478, 54.777218, 46.36312, 37.869293, 29.216341, 20.721802, 12.544483, 4.2080455, NaN, NaN, 100.21529, 94.85848, 87.95395, 78.07292, 67.9533, 57.952248, 48.90325, 39.496635, 29.851425, 20.563019, 11.631459, 5.2004952, 2.9377005, 1.9849374, NaN, NaN, 99.73912, 94.5807, 88.07298, 79.97772, 72.040886, 62.75439, 53.864365, 44.73581, 35.765614, 27.509512, 19.650028, 12.107817, 6.312033, 3.9301567, 3.3743815, NaN, NaN, 96.32663, 91.16813, 84.18411, 74.580696, 65.135574, 55.769394, 47.037823, 38.782177, 30.843742, 22.746222, 14.965948, 6.7090087, 1.7070467, NaN, NaN, 91.406204, 86.16822, 79.5015, 70.53283, 61.80189, 53.070576, 43.94199, 35.051147, 26.39808, 18.220995, 10.043581, 4.7241173, 2.42162, NaN, NaN, 96.52501, 92.00141, 86.36662, 77.63636, 68.90572, 60.49221, 52.157734, 43.66415, 35.17022, 27.15226, 19.213375, 11.036002, 5.1607943, 2.540715, 1.746745, NaN, NaN, 94.22353, 89.4618, 82.67614, 72.67581, 62.91311, 52.554615, 42.31467, 32.312366, 22.904993, 14.092629, 5.0417004, NaN, NaN, 92.27917, 87.2793, 81.009445, 72.596436, 64.26245, 55.13436, 45.847107, 36.797585, 28.065207, 19.253067, 9.805396, 3.5331728, 1.9452375, NaN, NaN, 91.644264, 86.80311, 80.53324, 71.96147, 63.548088, 54.737476, 46.085247, 37.6708, 29.335392, 20.602697, 11.3932705, 3.6919653, 1.4688544, NaN, NaN, 93.39023, 89.26338, 83.94598, 77.27918, 71.24714, 64.57993, 57.595013, 50.451096, 43.62445, 37.353264, 30.764341, 23.619488, 15.998035, 8.296904, 2.898, NaN, NaN, 90.612564, 85.69202, 79.025276, 69.18351, 59.261898, 49.498558, 40.68734, 31.95513, 23.540102, 15.362903, 7.661747, 4.24774, 2.7392068, 2.5010164, NaN, NaN, 95.53301, 92.19983, 87.04123, 78.549095, 69.50101, 60.61128, 52.03867, 44.02137, 36.003754, 28.700308, 21.872936, 15.601082, 9.0114565, 5.756263, 5.121097, NaN, NaN, 97.5964, 92.99346, 86.644424, 78.62847, 70.61221, 61.563778, 52.118057, 43.624474, 35.52746, 27.588896, 19.332466, 10.837521, 3.9301562, NaN, NaN, 99.2233, 93.74742, 86.68413, 77.47766, 68.66764, 59.301624, 50.570198, 41.917786, 33.66193, 25.643908, 18.101915, 10.321464, 4.8432136, 2.9377005, NaN, NaN, 101.127945, 95.41404, 88.27143, 78.35073, 68.42955, 58.50789, 49.06202, 39.774483, 30.96284, 22.70654, 14.608692, 7.3838716, 3.9698565, 2.3819232, NaN, NaN, 106.603645, 101.60412, 95.17598, 87.39845, 80.25556, 72.794945, 64.69908, 55.491623, 45.648712, 35.9641, 26.358412, 18.101925, 10.7978325, 3.8904612, NaN, NaN, 109.539856, 104.38168, 97.87427, 89.144485, 81.128624, 74.30299, 68.11211, 61.524162, 53.82473, 44.854923, 35.329037, 25.485155, 15.640799, 6.669319, 3.1758933, 2.0643363, NaN, NaN, 114.221825, 109.46054, 103.27072, 94.937965, 85.6525, 75.53324, 65.17536, 55.531353, 46.72038, 38.62347, 29.57361, 20.999687, 12.425406, 5.637179, 3.017101, 2.4216242, NaN, NaN, 118.66563, 113.78542, 107.23862, 98.78698, 89.73978, 80.09692, 69.97738, 60.09547, 50.68935, 43.06889, 36.757977, 30.56595, 22.944738, 14.8468895, 6.6296263, 1.6276528, NaN, NaN, 120.411415, 116.00737, 109.579666, 99.818695, 90.4144, 81.12872, 72.19978, 64.22294, 57.912678, 52.435688, 46.244137, 37.31368, 26.596617, 17.30804, 8.852691, 4.0889583, 2.1834345, NaN, NaN, 122.871346, 118.11027, 111.761986, 103.19149, 94.7, 85.73197, 76.525444, 66.92164, 57.396763, 48.18896, 39.457043, 31.201067, 22.150866, 13.020871, 5.9547696, 3.0171049, 1.8261477, NaN, NaN, 124.81548, 119.97509, 113.706215, 104.89773, 95.61269, 86.00978, 76.406425, 67.75507, 60.293987, 53.07076, 45.767895, 38.067856, 29.653048, 21.396673, 13.139966, 4.088962, NaN, NaN, 127.27536, 122.51438, 116.324936, 107.27848, 98.58875, 90.25579, 80.85104, 70.850586, 61.802128, 53.7058, 45.609154, 37.274036, 28.462257, 19.411926, 10.71847, 5.478399, 3.6919806, 3.2155998, NaN, NaN, 128.90205, 123.982414, 117.79301, 109.222755, 100.73151, 91.922455, 82.39873, 72.71581, 63.90556, 55.253674, 46.442665, 38.980793, 31.836195, 23.897457, 15.799628, 7.9396644, 3.8904738, 2.1437397, NaN, NaN, 129.93364, 125.17271, 118.74528, 108.984726, 98.74755, 87.79559, 77.55736, 68.03296, 59.34156, 52.316734, 44.815384, 36.480225, 27.430244, 18.0226, 9.090894, 2.7789185, NaN, NaN, 138.6221, 133.94072, 127.989655, 120.21334, 112.75415, 104.65983, 96.40646, 87.91467, 79.34316, 70.05696, 60.294083, 51.007015, 42.35458, 34.33686, 25.842497, 17.427172, 9.884843, 5.5975, 4.3271585, NaN, NaN, 134.21848, 129.53699, 123.34775, 115.3332, 107.873825, 100.09675, 91.76383, 82.875015, 74.462036, 65.33435, 55.650623, 46.36334, 37.79009, 29.534027, 21.59519, 13.73544, 6.986929, 4.5256515, 4.208065, NaN, NaN, 145.52507, 140.68515, 134.65494, 126.640816, 118.547035, 110.05616, 101.564926, 93.31143, 85.2957, 77.75587, 70.13638, 62.19912, 54.023415, 46.244286, 38.38548, 30.446985, 22.984518, 14.886641, 6.709047, 1.6276587, NaN, NaN, 147.8657, 143.1052, 136.75766, 128.90233, 122.71306, 116.444244, 109.461044, 101.366585, 92.71626, 83.827484, 75.17642, 66.445625, 57.873207, 49.53857, 41.679886, 33.423973, 24.135674, 15.243915, 7.78089, 4.605052, 3.9301803, NaN, NaN, 152.30882, 147.5484, 141.24068, 132.19531, 122.19732, 112.19885, 102.55701, 93.74801, 85.891014, 77.79562, 69.104614, 60.532307, 51.840572, 44.45826, 36.718452, 28.025707, 19.451677, 11.353653, 3.7316897, NaN, NaN, 157.62457, 152.46758, 146.19968, 138.66206, 131.67961, 124.062126, 116.285645, 108.508865, 100.7318, 93.0338, 85.65296, 78.351234, 71.12862, 64.14387, 57.000122, 49.697372, 41.20363, 32.8683, 25.485304, 17.943254, 10.440625, 5.7563043, 4.327168, 4.6050563, NaN, NaN, 162.7815, 158.02132, 151.83293, 143.97815, 136.20242, 128.18835, 120.412025, 112.79411, 104.77913, 96.84319, 88.58949, 79.93862, 71.44613, 63.588276, 56.127003, 48.98298, 41.36241, 33.662174, 26.914303, 20.324993, 12.782751, 5.6372123, 1.7467583, NaN, NaN, 174.68153, 169.44563, 163.01958, 154.84787, 147.07256, 138.26546, 129.53732, 120.88818, 112.47674, 104.38238, 96.20834, 87.87525, 79.621185, 71.36679, 63.588303, 56.127026, 48.1892, 40.5686, 33.26526, 25.72349, 17.784487, 10.083359, 5.557818, 4.208076, NaN, NaN, 181.34526, 176.42685, 169.76302, 161.03622, 152.30907, 143.26416, 134.45691, 126.04601, 117.71413, 109.54062, 101.9223, 94.62114, 86.84354, 78.510056, 69.938126, 61.842087, 54.30137, 47.157276, 39.933548, 32.550797, 25.247166, 17.466925, 9.845178, 3.33471, NaN, NaN, 184.55809, 179.71909, 173.68999, 165.36005, 156.79173, 148.06439, 139.65407, 131.08469, 122.91171, 114.42099, 106.00927, 97.8353, 89.74036, 81.96256, 74.025734, 65.929855, 57.833652, 50.134026, 42.83102, 35.845295, 28.899021, 21.754038, 14.370628, 8.0190935, 5.3990283, 4.9226494, NaN, NaN, 191.14217, 186.06532, 179.63979, 171.8654, 164.40805, 156.79176, 148.61981, 140.52687, 132.19557, 123.78459, 115.690674, 107.27901, 99.02572, 91.168915, 83.788, 76.168724, 68.628525, 60.532433, 52.912285, 45.450615, 37.8696, 30.248608, 22.547943, 15.323344, 7.9396996, 2.3025446, NaN, NaN, 193.44264, 188.84181, 182.73367, 174.7214, 166.78816, 158.21991, 149.6513, 141.16168, 132.83041, 124.1814, 115.37331, 107.12034, 98.78768, 90.93086, 82.83565, 74.263885, 66.08864, 57.833687, 49.65778, 41.87846, 34.257614, 26.47771, 19.173857, 11.552166, 3.8507946, NaN, NaN, 197.28983, 191.97517, 185.86711, 178.64825, 171.2705, 163.0991, 154.84807, 146.27931, 137.78957, 129.77554, 121.84055, 114.30204, 106.60453, 98.509926, 90.6531, 82.79597, 74.621056, 66.84269, 58.984642, 50.88816, 43.14858, 35.52778, 28.065474, 20.999847, 14.01337, 7.4236326, 4.724161, NaN, NaN, 214.77963, 209.70338, 202.56468, 194.31523, 186.3034, 177.89464, 169.72351, 161.55208, 153.22162, 145.12886, 136.87709, 128.78369, 120.76932, 112.75463, 104.898346, 96.88304, 89.10551, 81.089584, 73.07335, 65.215546, 57.397125, 49.697475, 42.076923, 34.85301, 28.105167, 21.754055, 15.085175, 8.336681, 3.017124, NaN, NaN, 255.42482, 250.30992, 243.41055, 232.94211, 222.83003, 212.95541, 204.38908, 196.53632, 188.80222, 180.82985, 172.26219, 163.57516, 154.76877, 145.96199, 137.39287, 128.70436, 120.015495, 111.56432, 103.35088, 95.25615, 87.31983, 79.62131, 72.39871, 64.858376, 57.476513, 50.173763, 42.870754, 35.88502, 29.13721, 22.62735, 15.879104, 9.130635, 5.7960157, 5.3990335, NaN, NaN, 333.56, 329.12085, 323.33395, 315.96136, 309.1435, 301.45328, 293.44562, 285.59625, 277.90515, 270.29306, 262.6014, 254.98874, 247.2172, 238.73161, 230.08705, 220.88693, 211.92435, 202.72342, 193.36343, 184.39966, 175.47514, 166.27258, 156.51425, 146.59676, 137.2342, 128.18863, 119.38071, 110.969185, 102.55732, 94.85937, 87.161125, 79.54196, 71.84314, 64.38215, 57.079647, 49.85626, 43.5852, 37.472717, 31.280664, 24.850258, 18.61813, 12.822475, 5.9151115, 1.945257, NaN, NaN, 392.2907, 385.5546, 378.81827, 371.0514, 363.522, 354.96194, 345.92593, 337.04807, 328.88324, 321.03522, 312.55267, 303.9112, 295.50723, 286.94434, 278.53967, 269.97607, 261.8879, 253.79941, 245.86922, 237.9387, 230.36479, 222.59232, 215.21611, 207.76033, 200.14565, 192.45134, 184.43945, 176.3479, 168.09738, 159.92586, 151.75401, 143.97856, 135.96477, 128.10938, 120.49172, 112.95315, 105.0175, 97.00219, 89.46275, 82.16113, 75.33547, 68.27147, 61.524723, 54.93651, 48.03056, 41.36253, 34.69428, 28.1052, 21.99225, 16.514257, 10.797935, 4.4462776, 1.2703749, NaN, NaN, 467.4038, 462.96753, 457.02594, 449.18277, 441.49777, 433.5748, 425.49304, 417.88638, 410.43793, 402.90997, 395.144, 387.53622, 379.84894, 371.92358, 363.91867, 355.9927, 348.06644, 340.37766, 332.6093, 324.7614, 316.83395, 309.30258, 301.8502, 294.55612, 287.02393, 279.9672, 273.1481, 266.48737, 259.74713, 253.00667, 246.10738, 239.12854, 232.14948, 225.17018, 218.03201, 210.73495, 203.19969, 195.5055, 187.89035, 180.2749, 172.73853, 165.43987, 158.0616, 150.9211, 143.701, 136.48067, 129.49811, 122.67402, 115.929054, 109.10451, 102.20038, 95.45474, 88.788246, 82.12154, 75.53397, 69.34306, 63.469463, 57.43694, 51.404236, 45.291977, 39.695526, 33.979847, 28.581556, 23.024343, 17.46698, 12.544619, 7.1457634, 2.937733, NaN, NaN, 501.94058, 497.58426, 491.64365, 482.5344, 473.50397, 464.63156, 456.07568, 447.51944, 438.72516, 429.9305, 421.45242, 412.89474, 404.3367, 396.01605, 387.61584, 379.21527, 370.81433, 362.49234, 354.09073, 346.00586, 338.11884, 330.19186, 322.2646, 314.17847, 306.25058, 298.48096, 290.7903, 283.0994, 275.3289, 267.32022, 259.46982, 251.61913, 243.53021, 235.20306, 226.79626, 218.46843, 210.21959, 201.89108, 193.7209, 185.47105, 177.57787, 169.96204, 162.66327, 155.36426, 148.06497, 140.76543, 133.62431, 126.086205, 118.54782, 110.77109, 103.15278, 95.931, 88.70896, 81.88351, 75.21657, 68.70815, 62.675777, 56.563847, 50.769253, 44.577587, 38.58419, 32.94786, 27.86709, 22.627415, 17.149427, 11.988872, 7.1457696, 3.096531, NaN, NaN, 500.59448, 495.68365, 489.1093, 480.55444, 471.91998, 463.60208, 455.52148, 447.51978, 439.5178, 431.11932, 422.95822, 414.71756, 406.47656, 398.23523, 390.07285, 381.5931, 372.87524, 364.3948, 356.23108, 348.14627, 340.2197, 332.2928, 324.4449, 316.51736, 308.431, 300.34433, 292.57446, 284.72504, 276.8753, 268.78738, 260.46124, 252.29338, 244.20448, 236.1946, 228.10507, 220.01523, 211.76643, 203.35867, 195.1092, 187.01807, 179.04561, 171.27116, 163.8931, 156.59412, 149.05684, 141.20192, 133.3467, 125.729225, 118.50823, 111.20763, 104.224205, 97.3199, 90.09791, 82.79629, 75.573784, 68.27165, 60.96926, 53.825367, 46.998745, 40.33066, 33.702053, 27.906805, 22.111395, 16.474606, 11.075845, 5.597545, 2.1040597, NaN, NaN, 501.22845, 496.7929, 490.69385, 482.37668, 474.13837, 465.89975, 457.26468, 449.0254, 440.78577, 432.46655, 423.98856, 415.35175, 406.5561, 398.15628, 389.7561, 381.6726, 373.66806, 365.4254, 357.10318, 348.54282, 340.18027, 331.53995, 322.97852, 314.33746, 305.8546, 297.21283, 288.72928, 280.0868, 271.8404, 263.75226, 256.06033, 248.606, 240.9928, 233.69655, 226.47934, 219.42052, 212.52008, 205.22282, 197.84598, 190.2309, 182.45686, 174.44455, 166.51126, 158.49834, 150.7231, 143.10628, 135.80653, 128.18915, 120.49213, 112.794815, 105.176575, 97.79613, 90.41542, 83.113815, 75.97069, 69.1448, 62.15993, 55.254204, 48.268864, 41.44205, 34.85317, 28.66101, 22.309887, 16.355528, 10.559787, 4.843278, 1.667371, NaN, NaN, 503.0505, 498.615, 492.6744, 484.991, 477.70337, 470.0194, 462.0975, 454.09604, 446.17352, 438.013, 429.77295, 421.6118, 413.4503, 405.12997, 396.8886, 388.64688, 380.3256, 372.00394, 363.84048, 355.5182, 346.91812, 338.4366, 329.95474, 321.7896, 313.38635, 305.37912, 297.29233, 289.0466, 280.95917, 272.8714, 264.86258, 256.8535, 249.00267, 241.15157, 233.37946, 225.52776, 217.75507, 209.90276, 202.44675, 195.06981, 187.97023, 180.75142, 173.6117, 166.55104, 159.56949, 152.42902, 145.12961, 137.75061, 130.13329, 122.277626, 114.818436, 107.59705, 99.978615, 93.07416, 86.56629, 79.97886, 73.1531, 66.723976, 60.612156, 54.341396, 48.070442, 41.719917, 35.845505, 29.4946, 23.540447, 17.90369, 12.425565, 6.709105, 2.7392468, NaN, NaN, 500.6747, 496.15994, 489.98166, 481.4268, 472.15863, 462.53354, 452.5515, 443.1632, 433.89334, 424.9796, 416.06546, 407.15097, 398.35495, 389.79626, 380.8806, 372.20236, 363.6426, 354.84473, 346.16537, 337.60455, 329.3208, 321.3935, 313.70367, 306.25143, 298.71964, 291.26685, 283.57593, 275.80542, 268.1932, 260.34283, 252.73006, 245.2756, 237.82088, 230.44519, 223.14856, 216.08961, 209.10974, 202.12962, 195.06995, 188.08936, 181.06888, 174.08781, 167.18584, 160.52165, 153.69856, 146.79591, 139.89304, 132.67252, 125.29306, 118.07204, 110.21591, 102.67692, 95.37574, 88.233025, 81.0107, 74.02623, 67.12089, 60.135944, 53.23014, 46.482864, 40.052902, 33.78151, 27.827475, 21.714489, 15.601319, 9.329176, 3.5332272, NaN, NaN, 498.06137, 493.38812, 487.36816, 479.28848, 471.05002, 462.81125, 454.9683, 447.28345, 439.2022, 431.43756, 423.59338, 415.59042, 407.5872, 399.58362, 391.42123, 383.41702, 375.25403, 367.32846, 359.32333, 351.15936, 343.1536, 335.06824, 327.06186, 318.9759, 311.12744, 303.43726, 295.90533, 287.81815, 279.88922, 272.19785, 264.2683, 256.4178, 248.72554, 241.03302, 233.65744, 226.3609, 218.82617, 211.37048, 204.15248, 196.8549, 189.2001, 181.58469, 174.12764, 166.90833, 159.37141, 152.07225, 145.16953, 138.58397, 132.15689, 125.65025, 119.38147, 112.47765, 105.9704, 99.78038, 93.43144, 86.923584, 80.57425, 74.30409, 68.27186, 62.3982, 56.405304, 50.451923, 44.339607, 38.147724, 32.431973, 26.636673, 20.761818, 14.966188, 9.329185, 3.7714238, NaN, NaN, 500.55676, 496.04196, 490.0221, 481.388, 472.67435, 463.485, 454.45367, 445.5804, 436.7068, 427.6743, 418.48294, 409.1327, 400.01974, 390.82718, 381.55493, 372.3615, 363.40546, 354.9246, 346.4434, 338.19965, 329.95554, 321.71112, 313.70422, 305.53842, 297.29303, 288.88873, 280.40482, 271.68265, 263.198, 254.79231, 246.70349, 238.77296, 230.76283, 222.83168, 214.6623, 206.65121, 198.63982, 190.54878, 182.61609, 174.84175, 166.9878, 159.13353, 151.19962, 143.42409, 135.96565, 128.34825, 120.65121, 112.795166, 105.01818, 97.79643, 90.97125, 83.90774, 77.00272, 70.335594, 63.43012, 56.762547, 50.174133, 43.664894, 37.23483, 30.96334, 24.890131, 19.174006, 13.934083, 7.9794626, 3.2156417, NaN, NaN, 499.0521, 494.14124, 487.72522, 479.48712, 471.72397, 463.56445, 455.32538, 447.00674, 438.5293, 429.9723, 421.49417, 413.0157, 404.93307, 396.7709, 388.7669, 380.6041, 372.44095, 364.436, 356.27225, 348.34592, 340.37967, 332.53204, 324.6048, 316.51874, 308.67017, 300.58347, 292.5757, 284.72626, 276.79718, 269.02643, 261.01746, 252.77026, 244.36415, 236.27492, 228.4233, 220.57137, 213.0364, 205.42186, 197.7277, 190.03326, 182.2592, 174.16753, 166.39287, 158.93526, 151.39804, 143.70186, 135.76735, 128.14993, 120.69094, 112.8349, 104.81984, 97.35999, 90.13797, 82.83633, 76.01064, 69.74034, 62.99359, 56.326, 49.81695, 43.307697, 36.996696, 30.80458, 24.53289, 18.816751, 13.179848, 7.4633913, 2.8583522, NaN, NaN, 499.40866, 494.577, 488.6363, 480.3982, 472.47665, 464.31717, 456.39502, 448.3933, 440.0744, 431.59668, 423.0394, 414.08554, 405.60675, 397.12762, 389.04437, 380.96082, 372.7977, 364.87204, 356.8668, 349.01978, 341.21207, 333.0474, 325.0409, 316.95483, 309.027, 301.25745, 293.329, 285.4003, 277.55054, 269.7798, 262.08804, 254.31671, 246.62437, 239.1697, 231.6354, 224.18018, 216.64536, 209.26889, 201.89217, 194.51517, 187.13791, 179.60173, 171.98593, 164.52853, 156.83284, 149.3749, 142.23404, 135.48969, 128.66574, 122.00029, 115.41397, 108.82744, 102.08198, 95.336296, 88.511024, 81.92363, 75.09791, 68.35134, 61.604546, 54.936905, 48.745335, 42.632954, 36.59978, 30.80459, 25.72374, 20.801546, 15.720448, 10.718618, 6.1930475, 2.5407603, NaN, NaN, 500.39896, 495.88416, 489.86426, 481.70544, 473.86316, 465.46606, 457.22705, 449.14615, 440.66882, 432.34958, 424.10925, 415.8686, 407.7861, 399.86176, 392.4126, 384.56693, 376.56247, 368.3199, 360.23553, 352.2301, 344.10547, 336.17868, 328.17233, 320.56204, 312.63434, 304.70636, 296.77805, 288.77017, 281.2377, 273.62567, 265.85477, 258.0836, 250.47069, 242.85753, 235.24406, 227.78896, 220.33359, 213.03656, 205.65997, 198.28311, 191.1043, 184.12355, 176.9839, 169.92336, 163.02122, 156.1982, 149.37495, 143.02754, 136.75928, 130.57018, 124.38089, 117.79464, 111.3669, 104.8596, 98.114, 91.68564, 85.018974, 78.3521, 71.764366, 65.17643, 58.548595, 51.880856, 45.054134, 38.941643, 32.749584, 26.795504, 21.158815, 15.363185, 9.884972, 5.1211896, 2.1040702, NaN, NaN, 500.20132, 495.44888, 489.11212, 480.39877, 471.3682, 462.25797, 453.46426, 444.74942, 435.95496, 427.3186, 418.60263, 410.04477, 401.56583, 393.00726, 384.3691, 375.6513, 367.09167, 358.76947, 350.5262, 342.2826, 334.27646, 326.27002, 318.184, 310.3355, 302.56598, 294.79614, 287.18463, 279.5728, 271.96072, 264.26904, 256.49777, 248.80553, 240.95436, 232.86499, 225.09253, 217.3198, 209.38812, 201.61478, 193.84114, 186.14655, 178.84831, 171.47047, 164.09238, 156.63469, 149.17671, 141.95651, 135.05344, 128.15013, 121.64335, 114.8983, 108.311745, 101.8837, 95.53481, 89.26509, 82.43961, 75.45516, 68.47048, 61.326805, 54.89728, 48.54694, 42.077324, 35.32966, 29.058096, 22.786343, 16.673183, 10.242259, 4.0493264, 0.8733909, NaN, NaN, 499.13226, 494.3006, 488.28064, 479.64645, 470.29898, 460.95105, 451.84036, 443.2839, 434.96475, 426.6453, 418.48395, 410.3223, 402.31882, 394.23578, 386.23166, 378.14798, 370.14325, 362.29672, 354.29135, 346.2857, 338.27972, 330.43198, 322.58395, 314.6563, 306.96625, 299.43445, 291.98163, 284.60788, 277.3131, 269.46304, 261.692, 253.84132, 246.06966, 238.37701, 230.60477, 222.51497, 214.42487, 206.49307, 198.56097, 190.7079, 182.85452, 175.00084, 167.2262, 159.37192, 151.59668, 143.97984, 136.36272, 128.904, 121.68308, 114.54126, 107.47854, 100.41558, 93.27302, 86.68577, 80.41577, 74.46307, 68.35145, 62.3984, 56.445175, 50.253635, 44.26037, 37.98908, 31.717594, 25.763477, 20.047361, 14.648662, 9.091027, 3.4538438, NaN, NaN, 498.37997, 493.46906, 487.29068, 479.60703, 472.0815, 464.31808, 456.31668, 448.47342, 440.7091, 433.10297, 425.49652, 417.73135, 410.12433, 402.51706, 394.83026, 387.2224, 379.45578, 371.68887, 364.00092, 356.2334, 348.5845, 341.05423, 333.52365, 326.0721, 318.62027, 310.93033, 303.16083, 295.4703, 287.70023, 279.69196, 271.9213, 264.1503, 256.2997, 248.29025, 240.67699, 233.06345, 225.3703, 217.7562, 210.6177, 203.32034, 196.22102, 188.92313, 181.86298, 174.6439, 167.50392, 160.3637, 153.22322, 146.32051, 139.65562, 132.91116, 125.92842, 119.10416, 111.96224, 104.89944, 98.15383, 91.487366, 84.66196, 77.677574, 71.01045, 64.6606, 58.350246, 52.079384, 46.046474, 40.01339, 33.741966, 27.708517, 22.230627, 16.831982, 11.988959, 6.7488384, 2.5407653, NaN, NaN, 500.28116, 495.52872, 489.4296, 481.5084, 473.98294, 466.14038, 458.21826, 449.97894, 441.66006, 433.34085, 425.4175, 417.49384, 409.8076, 402.0418, 394.19647, 386.2716, 378.50494, 370.81723, 363.2085, 355.52023, 347.75238, 340.06354, 332.29514, 324.52643, 316.8367, 309.1467, 301.61496, 294.08298, 286.62997, 278.93884, 271.4853, 264.19006, 256.8153, 249.59886, 242.6201, 235.6411, 228.89978, 222.23756, 215.25786, 208.1193, 201.25809, 194.19835, 187.05905, 179.99883, 172.93835, 165.95697, 158.73735, 151.59682, 144.13864, 137.07695, 129.85631, 122.55605, 115.41425, 108.27221, 100.89183, 93.908, 86.923935, 80.41584, 73.98691, 67.95464, 61.72376, 55.77051, 50.13461, 44.49855, 38.782955, 33.305355, 27.748224, 22.508505, 17.189259, 11.711083, 5.835776, 2.2628717, NaN, NaN, 497.90527, 492.99435, 486.4991, 478.02325, 470.0224, 461.86276, 454.0197, 446.09714, 437.93655, 429.93414, 421.77292, 413.53214, 405.29105, 397.04962, 388.7286, 380.4865, 372.24408, 364.15985, 356.0753, 347.99042, 340.02414, 332.01788, 323.93207, 316.0045, 307.83878, 299.98987, 292.14066, 284.529, 276.6792, 269.22556, 261.85095, 254.4761, 247.33888, 240.20142, 232.74648, 225.37056, 217.75644, 210.53864, 203.16193, 195.70564, 188.28873, 180.99055, 173.93011, 166.94878, 160.04652, 153.06471, 146.00331, 138.94167, 131.80043, 125.61116, 120.45329, 115.45401, 110.53395, 105.534424, 100.534775, 95.376274, 90.13828, 84.900154, 79.74126, 75.05846, 70.534294, 66.01003, 61.7238, 57.199345, 52.51603, 47.515083, 42.593395, 37.59221, 32.511513, 27.510077, 22.429129, 17.586233, 12.981406, 7.661908, 3.1362562, NaN, NaN, 500.47983, 495.7274, 489.54904, 481.86548, 474.02316, 465.94293, 457.94156, 449.9399, 441.70026, 433.38104, 425.0615, 416.7416, 408.4214, 400.18005, 392.17618, 384.33044, 376.48447, 368.47964, 360.31598, 352.6276, 345.1371, 337.60666, 329.83813, 322.54498, 314.93445, 307.32364, 300.0297, 292.33905, 284.72742, 276.95688, 269.26538, 261.4943, 253.6436, 246.03053, 238.33786, 230.64491, 223.03098, 215.57541, 207.96092, 200.42548, 193.08806, 185.6314, 178.33311, 170.87592, 163.41844, 155.88136, 148.18532, 140.96506, 133.74455, 126.52377, 119.54081, 112.63696, 105.57417, 98.59049, 91.765305, 85.098625, 78.431725, 72.08209, 65.73227, 59.382244, 53.389233, 47.197586, 40.926373, 34.258038, 28.065815, 21.952797, 15.839597, 9.567422, 3.8508418, NaN, NaN, 500.5592, 495.80676, 489.54922, 481.07352, 472.75586, 464.67557, 456.1196, 447.48407, 438.61047, 429.89496, 421.09982, 412.2251, 403.03302, 394.1575, 385.83636, 377.43564, 368.71753, 360.3161, 352.07288, 343.75003, 335.50613, 327.2619, 318.8588, 310.77243, 302.6065, 294.7574, 286.98724, 279.2961, 271.76328, 264.30945, 256.61746, 248.8459, 241.54987, 234.17427, 227.03635, 219.97748, 212.91838, 205.70038, 198.72011, 191.50163, 184.24323, 176.86557, 169.56697, 162.03012, 154.731, 147.51097, 140.13199, 133.07014, 125.690636, 118.786995, 111.96248, 105.13773, 98.2334, 91.328835, 84.7415, 78.23333, 71.24872, 64.184494, 57.358154, 50.61097, 43.546036, 36.480854, 29.891758, 23.38184, 17.0305, 10.75836, 4.803618, 1.4688869, NaN, NaN, 497.78714, 492.9554, 486.61856, 477.9051, 469.03278, 459.764, 450.97015, 442.0175, 433.3021, 424.58636, 415.79102, 407.15378, 398.83316, 390.82922, 382.82495, 374.97888, 367.37027, 359.99918, 352.7071, 345.33548, 338.12213, 330.51218, 322.9812, 315.3707, 307.3635, 299.67313, 292.06174, 284.5294, 277.07602, 269.38452, 261.9306, 254.39714, 246.78409, 239.25006, 231.79506, 224.26048, 216.88426, 209.5871, 202.13103, 194.91266, 187.45605, 179.99918, 172.78003, 165.4813, 158.26163, 150.64502, 143.34549, 135.88701, 128.50761, 121.52472, 114.54158, 107.47884, 100.574585, 93.27328, 86.44791, 79.86042, 73.828316, 68.113525, 62.557323, 57.080353, 51.603233, 46.205353, 40.64856, 34.77407, 29.137579, 23.659714, 18.102308, 12.465358, 6.431267, 2.4613729, NaN, NaN, 499.64868, 494.6586, 488.24258, 479.1331, 469.6271, 460.83368, 452.1983, 443.8003, 435.24344, 427.0032, 418.9211, 410.83868, 402.83517, 394.59363, 386.27252, 377.79254, 369.47073, 361.06934, 352.6676, 344.42404, 335.70453, 327.4603, 319.21576, 311.12943, 303.43918, 295.74866, 288.05783, 280.28745, 272.51675, 264.98367, 257.45032, 249.99597, 242.38275, 234.92787, 227.3934, 219.93797, 212.72023, 205.18495, 197.72871, 190.58951, 183.48973, 176.42937, 169.28943, 162.0699, 154.77078, 147.4714, 140.2511, 133.18925, 126.206505, 119.38223, 112.47837, 105.17749, 97.79698, 90.01939, 82.162125, 74.78079, 67.47856, 60.25545, 52.873325, 46.046604, 39.735657, 33.464207, 27.271955, 21.397081, 15.680826, 9.805619, 4.48603, 1.3894888, NaN, NaN, 497.86667, 492.95572, 486.53967, 478.22223, 470.459, 462.22015, 454.0602, 445.8207, 437.42242, 429.34073, 421.33795, 413.2556, 405.33145, 397.09003, 389.08597, 381.08163, 373.394, 365.7061, 357.93863, 350.17087, 342.3632, 334.7534, 326.9055, 318.978, 311.05023, 303.12213, 295.19373, 287.10645, 279.09814, 270.85165, 262.7634, 254.67485, 246.9825, 239.21056, 231.67624, 224.14166, 216.21022, 208.67506, 201.21895, 193.76257, 186.42491, 179.28532, 172.14548, 165.16406, 158.26173, 151.35918, 144.53574, 137.55338, 130.65013, 123.74665, 116.60487, 109.30414, 102.16186, 95.49551, 88.670204, 82.08278, 75.49515, 68.19294, 60.890472, 53.825886, 47.118267, 40.52951, 33.781765, 27.113184, 21.079521, 15.045681, 8.297095, 3.0568638, NaN, NaN, 499.56976, 494.7381, 488.40128, 479.52942, 470.81564, 462.10147, 453.70386, 445.54355, 437.5414, 429.61816, 421.53616, 413.7708, 405.76743, 397.68448, 389.60123, 381.67615, 373.59225, 365.66656, 357.58206, 349.5765, 341.61026, 333.68335, 326.0732, 318.22498, 310.535, 302.84473, 295.0749, 287.38403, 279.8515, 272.1601, 264.70627, 257.1729, 249.71855, 242.58115, 235.44351, 228.14699, 220.92953, 213.7118, 206.41452, 199.27562, 192.25546, 185.19539, 178.29375, 171.2332, 164.72775, 158.14278, 151.63692, 145.13086, 138.54526, 132.11812, 125.690796, 119.02521, 111.88326, 104.74107, 97.757355, 91.01149, 84.50351, 78.3128, 72.04253, 65.61331, 58.826706, 52.23832, 46.04663, 39.93414, 34.059628, 28.264332, 22.548265, 16.832039, 11.353839, 5.557902, 1.9055834, NaN, NaN, 500.04517, 495.53033, 489.5896, 481.2723, 472.87546, 464.00293, 455.60538, 447.36594, 438.88846, 430.80682, 422.72485, 414.4841, 406.4015, 398.39783, 390.47308, 382.46878, 374.6227, 366.6178, 358.69183, 350.84485, 343.03717, 335.26886, 327.65878, 319.96915, 312.12067, 304.2719, 296.34357, 288.4149, 280.32733, 272.31876, 264.072, 255.66628, 247.18092, 238.85382, 230.36777, 222.04, 213.47394, 205.06615, 196.896, 188.88417, 181.07036, 173.37524, 165.83852, 158.53952, 151.31961, 143.8614, 136.1649, 128.54745, 120.77102, 113.153, 105.85213, 98.551, 91.40834, 84.42417, 77.677864, 70.93134, 64.343346, 57.675755, 50.84919, 44.339928, 37.87015, 31.598642, 26.200224, 21.039839, 15.720537, 9.845326, 3.8905485, NaN, NaN, 500.79782, 496.2038, 490.10464, 481.23288, 472.43994, 463.9635, 455.40747, 447.32648, 439.64133, 432.0351, 424.34937, 416.58408, 408.66006, 400.65646, 392.65256, 384.64835, 376.3268, 368.32196, 360.31683, 352.07358, 344.06778, 336.06168, 328.2138, 320.36566, 312.43793, 304.50986, 296.5815, 288.57358, 280.5653, 272.55676, 264.30997, 256.30078, 248.29126, 240.36075, 232.03337, 224.02292, 216.09146, 208.31833, 200.86221, 193.4058, 186.14746, 179.08717, 171.94731, 164.72787, 157.50818, 150.44691, 143.06802, 135.68887, 128.30945, 120.771065, 113.2324, 105.53474, 97.75742, 90.53537, 83.392426, 76.16987, 69.1058, 62.279613, 55.691334, 49.02346, 42.672905, 36.163383, 29.971203, 24.01701, 17.98325, 12.028706, 6.2327843, 2.3422787, NaN, NaN, 498.58038, 493.74866, 487.57025, 479.17365, 470.61826, 462.0625, 453.5064, 444.87073, 436.71008, 428.5491, 420.5463, 412.46393, 404.38123, 396.0605, 387.8979, 379.735, 371.17548, 362.53635, 353.8176, 345.33627, 336.8546, 328.2933, 319.89023, 311.56607, 303.40012, 295.31317, 287.30518, 279.37613, 271.6847, 263.91367, 256.53885, 249.24307, 241.86774, 234.57144, 227.19557, 219.97806, 212.2844, 204.66977, 197.05486, 189.59831, 182.06216, 174.20842, 166.51305, 158.97604, 151.6768, 144.61533, 137.39493, 130.17426, 122.79464, 115.65282, 108.19331, 100.65418, 92.87668, 85.257614, 78.43196, 72.00294, 65.41497, 59.22367, 53.111565, 47.316803, 42.07756, 36.52064, 31.201736, 25.962084, 20.722296, 15.402979, 9.924733, 4.684534, 1.5085905, NaN, NaN, 501.66983, 497.31342, 491.37274, 483.1347, 474.7379, 466.26157, 457.86407, 449.38702, 440.90964, 432.19418, 423.55762, 415.1584, 406.3626, 397.88345, 389.40393, 381.16183, 372.9194, 364.51813, 355.95798, 347.4767, 339.27258, 331.187, 323.1804, 315.0942, 307.16626, 299.1587, 291.23013, 283.14267, 274.97562, 266.7289, 258.7991, 250.78967, 242.46272, 234.37334, 226.6009, 218.74886, 211.05513, 203.36113, 195.66684, 187.89293, 180.19806, 172.34424, 164.25209, 156.31831, 148.78094, 141.16396, 133.70538, 126.24653, 118.86676, 111.64544, 104.66194, 97.99565, 91.40851, 85.05926, 78.86855, 72.43954, 66.0897, 60.05717, 54.42136, 48.54725, 42.71266, 37.155754, 31.519312, 25.962103, 20.484135, 15.561778, 10.004136, 4.6845374, 1.5879908, NaN, NaN, 497.78897, 493.11566, 486.9372, 478.699, 470.6189, 462.45923, 454.45773, 446.29742, 437.97836, 429.89667, 421.9731, 413.8908, 406.0459, 398.35916, 390.51364, 382.66785, 374.901, 367.13385, 359.28717, 351.51944, 343.7118, 336.18127, 328.57123, 320.96088, 313.35025, 305.81863, 298.4453, 290.99243, 283.69788, 276.32376, 269.0287, 261.73334, 254.35843, 246.74535, 239.29059, 231.91489, 224.85616, 217.47993, 210.26207, 203.12329, 195.8256, 188.60698, 181.3881, 174.40698, 167.10828, 159.88866, 152.82745, 145.84535, 139.02171, 132.27719, 125.61179, 118.86683, 112.28036, 106.16982, 99.74166, 93.23394, 86.646645, 80.138504, 73.31267, 66.80411, 60.49378, 54.699215, 48.90449, 43.34775, 38.26717, 33.02769, 28.105633, 23.501019, 18.81691, 13.815115, 8.575009, 3.6523626, NaN, NaN, 499.13574, 494.30405, 488.28406, 480.0459, 471.8074, 463.17245, 454.53717, 446.13922, 437.58243, 429.50073, 421.33945, 412.8609, 404.382, 396.3782, 388.29486, 380.0527, 371.96872, 363.9637, 356.03763, 348.11124, 340.66016, 333.12952, 325.3608, 317.82962, 310.13962, 302.37003, 294.6794, 287.2264, 279.69382, 272.08167, 264.46924, 257.09445, 249.71936, 242.34402, 234.96841, 227.51324, 220.1371, 212.91934, 205.54268, 198.24507, 191.0662, 184.00607, 177.02502, 169.96442, 162.50687, 155.28708, 148.14638, 140.92607, 133.54683, 126.08796, 119.10495, 112.1217, 105.05885, 98.15448, 91.01179, 83.47201, 76.56692, 69.42347, 62.756027, 56.088367, 49.618942, 43.189007, 36.600098, 30.24914, 24.215548, 18.181778, 12.386015, 7.2252665, 3.0171752, NaN, NaN, 499.136, 494.3835, 488.36353, 480.36298, 472.75824, 464.99478, 457.23102, 449.46698, 442.01956, 434.73032, 427.20312, 419.67566, 412.22717, 404.69916, 397.5671, 390.19705, 382.906, 375.45618, 368.24384, 360.63495, 352.58984, 344.66333, 336.65723, 328.49228, 320.2477, 311.76498, 303.28192, 295.03635, 286.94904, 278.7821, 270.61487, 262.4473, 254.27937, 246.26976, 238.49776, 230.88408, 223.42874, 216.2904, 209.15182, 202.01299, 194.55661, 187.41727, 180.51567, 173.69316, 166.94978, 160.04749, 153.30365, 146.63893, 139.8153, 133.15015, 126.802185, 120.29531, 113.47081, 106.8048, 100.05921, 93.23403, 86.7261, 80.6148, 74.8208, 69.18538, 63.62919, 57.83471, 51.643166, 44.975143, 38.386288, 32.273544, 26.636957, 20.76204, 15.283924, 9.805662, 4.724244, 1.5482937, NaN, NaN, 500.95795, 496.36392, 490.26477, 481.78903, 473.23373, 464.28198, 455.09216, 446.21884, 437.2659, 428.3918, 419.5966, 410.88022, 402.08426, 393.4464, 384.88742, 376.64514, 368.48175, 360.3973, 352.3918, 344.38602, 336.34027, 328.4924, 320.80276, 313.19214, 305.81906, 298.44574, 290.99286, 283.77756, 276.32416, 269.10834, 261.8923, 254.67598, 247.61803, 240.48053, 233.26347, 226.12547, 218.98723, 212.166, 205.02727, 197.80898, 190.7094, 183.33194, 176.27153, 169.13155, 162.07066, 154.93019, 147.55144, 140.25177, 132.79314, 125.81035, 118.35119, 111.05048, 103.74951, 95.81338, 88.4325, 81.05135, 73.98743, 67.55825, 61.525753, 55.49308, 49.182392, 42.9112, 37.116135, 31.241516, 25.6049, 19.968126, 14.410593, 8.455926, 3.1362762, NaN, NaN, 500.1264, 495.2947, 489.27475, 480.64053, 471.6099, 462.8165, 454.18118, 445.86243, 437.54333, 429.38235, 421.45877, 413.3764, 405.29373, 397.21075, 389.36517, 381.44006, 373.4354, 365.43042, 357.26657, 349.34024, 341.29468, 333.20917, 325.12335, 317.19577, 309.26788, 301.3397, 293.56976, 285.8788, 278.1083, 270.4961, 262.8043, 255.11221, 247.02332, 239.09271, 231.0825, 222.91335, 214.50592, 206.41544, 198.2453, 190.07484, 182.10237, 174.24861, 166.5532, 158.77818, 151.47891, 144.17937, 136.95892, 129.57953, 122.43792, 115.216705, 108.39204, 101.72585, 95.29755, 89.02776, 82.59906, 76.011406, 69.50292, 63.0736, 56.96159, 51.16692, 45.491158, 39.378624, 33.107132, 26.75606, 20.404789, 14.291506, 7.6222606, 2.699583, NaN, NaN, 499.80975, 495.13647, 488.79965, 480.48227, 472.00613, 463.37122, 454.89438, 446.17947, 437.8604, 429.7787, 421.6174, 413.4558, 405.6901, 398.08258, 390.55405, 383.02524, 375.49615, 367.88754, 360.19937, 352.74872, 345.13928, 337.52954, 329.99878, 322.07138, 314.14368, 306.61206, 299.39734, 291.94446, 284.57065, 277.19653, 269.66357, 261.97174, 254.35893, 246.58722, 238.89453, 231.20155, 223.34966, 215.89404, 208.43816, 200.90268, 193.32727, 185.7119, 178.33426, 170.877, 163.49883, 155.80302, 148.10692, 140.33119, 132.71387, 125.09626, 117.55772, 110.018906, 102.717896, 95.41662, 88.03572, 80.89267, 74.06685, 67.637665, 61.049534, 54.38181, 48.26954, 42.23647, 36.44138, 30.40796, 24.533146, 18.89634, 13.179984, 7.2252774, 2.858382, NaN, NaN, 501.8694, 497.43378, 491.57227, 483.8095, 476.2841, 468.59998, 460.6779, 452.9932, 444.99127, 436.98907, 428.98654, 420.82523, 412.6636, 404.50165, 396.02237, 387.78052, 379.45905, 371.13727, 362.8944, 354.80975, 346.72476, 338.71875, 330.79166, 322.94357, 315.17444, 307.40503, 299.7146, 292.10318, 284.4915, 276.8795, 269.26724, 261.57538, 254.04185, 246.42874, 238.97395, 231.67752, 224.22221, 217.16321, 209.70737, 202.48921, 195.15182, 187.85385, 180.5556, 173.17776, 165.48232, 158.0246, 150.64595, 143.18768, 135.57047, 127.714905, 119.70034, 111.76482, 103.82899, 96.051575, 88.51196, 81.051445, 73.59065, 66.68521, 60.097046, 53.508667, 47.237602, 41.2045, 34.93306, 28.661427, 22.548384, 16.514553, 10.798127, 5.002145, 1.6673951, NaN, NaN, 499.96872, 495.45386, 489.5131, 481.43338, 473.59103, 465.51068, 457.43005, 449.4283, 441.34702, 433.34467, 425.5797, 417.89368, 410.12814, 402.44153, 394.83392, 387.0675, 379.22153, 371.37527, 363.60797, 355.6026, 347.63654, 339.47202, 331.30713, 322.82486, 314.4215, 306.25565, 298.16876, 290.16083, 281.99402, 273.82687, 265.6594, 257.4916, 249.5614, 241.47227, 233.70007, 225.76895, 217.91684, 209.9851, 202.37036, 194.83466, 187.61598, 180.07973, 172.70187, 165.32375, 158.02469, 150.88406, 143.66385, 136.36403, 128.8259, 121.44619, 113.98686, 106.44791, 98.67059, 91.051704, 83.750015, 76.84491, 69.8602, 63.11338, 56.604473, 50.174736, 44.022644, 37.433743, 31.082794, 24.89043, 18.777271, 12.981511, 6.709202, 2.3422909, NaN, NaN, 500.52344, 495.92935, 489.9094, 482.14658, 474.54187, 466.85767, 459.09396, 451.25073, 443.56567, 435.72186, 427.7985, 419.79562, 411.79242, 403.70966, 395.78506, 387.78094, 379.7765, 371.93027, 363.84595, 355.7613, 347.59708, 339.43253, 331.5055, 323.49887, 315.1748, 307.08826, 299.00137, 291.31064, 283.6196, 275.849, 268.15738, 260.2276, 252.05959, 244.12917, 236.27774, 228.42603, 220.41539, 212.3251, 204.39316, 196.69887, 189.28194, 181.66643, 174.20929, 166.8312, 159.45287, 151.83624, 143.8226, 136.0467, 127.9531, 120.335304, 112.717224, 105.41629, 98.27383, 91.52794, 85.178665, 78.670456, 72.24142, 66.20904, 60.335243, 54.14376, 47.872707, 41.998386, 36.123894, 30.40801, 24.453794, 18.658192, 13.021215, 6.748904, 2.7789874, NaN, NaN, 498.5435, 493.63254, 487.1372, 478.58212, 470.42276, 462.0254, 453.2316, 444.35815, 435.64282, 426.92712, 418.44876, 409.73233, 400.93628, 391.74362, 383.2638, 374.62512, 366.22388, 357.74304, 349.18256, 340.78027, 332.13983, 323.57828, 314.85785, 306.45413, 297.89154, 289.2493, 280.76526, 272.28088, 263.79617, 255.62828, 247.5394, 239.6088, 231.6779, 223.74669, 215.9738, 208.27995, 200.42715, 192.73273, 185.11732, 177.81897, 170.71869, 163.65784, 156.59674, 149.45605, 142.23578, 134.7772, 127.15965, 119.85924, 112.39985, 105.09891, 98.27388, 91.369255, 84.38503, 77.24184, 70.25713, 63.351566, 56.44577, 49.61912, 42.95101, 36.759, 31.162212, 25.128626, 19.65061, 14.331238, 8.455949, 3.2950826, NaN, NaN, 500.24673, 495.41504, 489.31586, 480.76083, 471.88858, 462.93674, 454.3014, 446.06186, 437.9804, 429.89868, 421.9751, 414.13046, 406.20627, 398.44028, 390.8325, 383.2244, 375.61606, 368.16592, 360.71555, 353.34415, 345.93286, 338.56094, 330.95093, 323.1821, 315.25443, 307.56427, 299.87384, 292.02454, 284.17496, 276.40436, 268.71274, 261.10016, 253.40799, 245.71553, 238.1814, 230.7263, 223.19162, 215.57735, 208.20076, 200.58592, 193.05014, 185.67274, 178.3744, 171.0758, 163.6976, 156.16046, 148.86108, 141.48209, 134.18217, 127.0407, 119.89899, 112.75702, 105.535446, 98.313614, 91.32963, 84.90098, 78.71023, 72.91615, 67.59816, 62.438786, 57.120518, 51.484596, 45.9279, 39.97413, 33.782024, 28.304237, 22.905695, 17.189436, 11.314225, 5.041855, 1.9452972, NaN, NaN, 496.99945, 492.08847, 485.5931, 477.19638, 468.72006, 460.08496, 451.4495, 443.05136, 434.8906, 426.7295, 418.96426, 411.1195, 403.3537, 395.74606, 387.97968, 380.21298, 372.20825, 364.2032, 356.03928, 348.11285, 340.22577, 332.0609, 323.975, 315.96808, 307.96082, 300.429, 292.73828, 285.12656, 277.6732, 269.9023, 262.13116, 254.51834, 247.22244, 239.76767, 232.31264, 224.61938, 216.84653, 208.91473, 201.45857, 194.08147, 186.66443, 179.44545, 172.46422, 165.40343, 158.26303, 150.56702, 142.95004, 135.33278, 127.71525, 120.09743, 112.479324, 105.3371, 98.51207, 92.00427, 85.57564, 78.98806, 72.95588, 66.76476, 60.49409, 54.54074, 48.626907, 42.99075, 38.068905, 33.067554, 27.589746, 21.794224, 15.998536, 10.52027, 4.4066696, 1.2307011, NaN, NaN, 500.92044, 496.16797, 490.0688, 481.43457, 472.64157, 463.76898, 454.97522, 446.33954, 437.9412, 429.62173, 421.22272, 413.21954, 405.29532, 397.13306, 389.20822, 381.3623, 373.43686, 365.35257, 357.50577, 349.65866, 341.9698, 334.35992, 326.67047, 319.06003, 311.21146, 303.67972, 295.98914, 288.45685, 280.7657, 273.07425, 265.30322, 257.6905, 249.99818, 242.3056, 234.61272, 226.99886, 219.3054, 211.61166, 203.99695, 196.22331, 188.56837, 180.79414, 172.94029, 165.0068, 157.62839, 150.32904, 142.95009, 135.57088, 128.1914, 120.49425, 113.272934, 106.36881, 99.543816, 92.63923, 85.813774, 79.226204, 72.79716, 66.60604, 60.33536, 54.143867, 47.872803, 41.522163, 35.250713, 29.296627, 23.818714, 18.499443, 12.862451, 7.1459055, 3.0171905, NaN, NaN, 499.01962, 494.2671, 488.08862, 478.82062, 468.8392, 459.4515, 449.94452, 440.91248, 431.9989, 423.08493, 414.28943, 405.49356, 396.8162, 388.01956, 379.22256, 370.90076, 362.34082, 354.1372, 346.17108, 338.20462, 330.2775, 322.58792, 314.97733, 307.36642, 299.75528, 292.3024, 284.92853, 277.39584, 269.62497, 261.7745, 254.00305, 246.23131, 238.14203, 230.13174, 222.20045, 214.11024, 205.86105, 197.69087, 189.679, 181.66682, 173.89235, 166.1969, 158.97719, 151.91592, 145.01309, 138.58612, 132.07959, 125.41415, 119.06591, 112.4794, 105.65461, 98.5915, 91.60751, 84.78202, 78.432526, 71.84471, 65.653564, 59.700363, 53.746986, 48.269726, 42.99078, 37.51323, 32.2737, 26.716476, 21.159101, 16.077942, 10.758466, 5.5976486, 2.3422973, NaN, NaN, 500.08914, 495.33664, 489.15823, 480.76163, 473.07764, 465.631, 458.0257, 450.34085, 442.735, 435.1288, 427.52234, 419.91562, 412.22937, 404.54282, 396.93524, 389.08963, 381.40222, 373.87305, 366.42285, 358.81387, 351.36313, 343.9914, 336.46085, 329.16785, 321.4782, 313.94684, 306.49448, 299.04184, 291.58896, 284.13577, 276.8409, 269.5458, 262.25043, 254.8755, 247.6589, 240.44206, 233.22498, 226.24556, 219.1866, 211.81012, 204.711, 197.6513, 190.4327, 183.21385, 175.83607, 168.77538, 161.79378, 154.89128, 148.0679, 141.16493, 134.0237, 127.04092, 120.05789, 113.15399, 106.48793, 100.13911, 93.869446, 87.75832, 81.726395, 76.011765, 70.61447, 65.21703, 59.50195, 53.7867, 48.150677, 42.673264, 37.195705, 31.638613, 26.001978, 20.76215, 15.760372, 10.679075, 5.5976515, 2.0247002, NaN, NaN, 499.1389, 494.38635, 488.1287, 479.9697, 471.49347, 463.17538, 454.6985, 446.30048, 437.9021, 429.6619, 421.42133, 413.1012, 404.7015, 396.30145, 388.05954, 380.13434, 372.12958, 364.20377, 356.67395, 348.98535, 341.29645, 333.36945, 325.60068, 317.59378, 309.983, 302.4512, 294.76056, 287.2282, 279.93347, 272.47986, 265.1846, 257.57187, 249.64163, 241.71109, 233.85956, 225.9284, 218.39354, 210.8584, 203.16432, 195.54929, 188.33061, 181.19102, 174.3685, 167.62509, 160.9608, 154.2963, 147.47289, 140.5699, 133.42865, 126.68389, 119.85956, 113.035, 106.60702, 100.099464, 93.512344, 86.92501, 79.86125, 73.35285, 67.003, 60.89107, 55.017105, 49.142967, 43.824345, 38.50559, 33.345467, 28.105824, 22.866047, 17.70553, 12.544884, 7.3047094, 2.937795, NaN, NaN, 498.86252, 494.11, 488.08994, 479.85168, 471.61313, 463.37424, 455.29346, 446.97467, 438.7348, 430.57382, 422.41254, 414.33014, 406.3267, 398.4814, 390.47736, 382.71072, 374.7853, 366.8596, 358.93353, 350.7694, 343.1202, 335.3518, 327.5038, 319.25916, 311.41058, 303.40314, 295.6332, 287.78372, 279.93393, 272.16315, 264.39206, 256.69998, 249.16623, 241.47359, 233.78065, 226.24606, 218.71118, 211.17604, 203.9579, 196.97748, 189.99681, 182.53995, 174.92413, 167.46672, 160.00902, 152.78908, 145.80693, 138.90387, 132.318, 125.96995, 119.383644, 113.35263, 107.321434, 101.13134, 94.623604, 87.95693, 81.05193, 74.62293, 68.669975, 63.193096, 57.795452, 52.159527, 46.126534, 40.4109, 34.93327, 29.693659, 24.612696, 19.928574, 15.323736, 10.480607, 5.5579643, 2.0644045, NaN, NaN, 497.71515, 492.9626, 486.78406, 479.02106, 471.8123, 464.3656, 456.68094, 449.2337, 441.94467, 434.89307, 427.762, 420.4722, 413.18213, 405.8918, 398.68048, 391.3104, 383.8608, 376.80722, 369.59485, 362.22372, 355.1694, 347.87704, 340.66367, 333.3708, 326.15692, 318.9428, 311.887, 304.67236, 297.4575, 290.32166, 283.02698, 275.89066, 268.59546, 261.61722, 254.79735, 248.05655, 241.39485, 234.89154, 228.54666, 221.88431, 215.34073, 208.83661, 202.33228, 195.82773, 189.08499, 182.34204, 175.6782, 169.25215, 162.74657, 156.39944, 149.89345, 143.54594, 137.19823, 130.61227, 124.26417, 117.8365, 111.80543, 105.77418, 99.66338, 94.028595, 88.03651, 82.004555, 76.21053, 70.65448, 65.336395, 59.780037, 54.144154, 48.34935, 42.71315, 37.6325, 32.472332, 27.391428, 22.469181, 17.62621, 12.703727, 7.463535, 3.0172064, NaN, NaN, 499.53815, 494.94403, 488.92398, 480.6065, 472.13028, 463.7329, 455.0183, 446.38257, 437.74646, 429.03076, 420.47318, 411.75674, 403.19846, 394.4813, 386.00153, 377.36288, 368.4861, 359.7675, 351.0485, 342.72546, 334.56067, 326.63333, 318.94357, 311.33276, 303.80096, 296.3482, 288.4987, 280.8075, 273.43317, 266.0586, 258.28723, 250.35698, 241.79196, 233.54382, 225.61261, 217.83974, 210.2252, 202.76903, 195.47124, 188.17317, 181.03352, 173.65562, 166.3568, 159.37506, 152.71046, 145.80762, 138.26974, 130.5729, 123.03449, 115.73386, 108.829765, 102.16352, 96.052605, 89.70341, 83.27465, 76.92506, 70.57527, 64.701546, 58.907024, 53.42986, 48.309772, 43.229248, 37.513508, 32.11516, 26.557892, 21.159258, 15.601691, 10.043973, 4.8831, 1.7865134, NaN, NaN, 498.78644, 494.1131, 488.0138, 479.77548, 471.53687, 463.2979, 454.90018, 446.5021, 438.18292, 429.70496, 421.54358, 413.38187, 405.21982, 397.05746, 388.81555, 380.81107, 372.727, 364.80115, 357.2713, 349.82043, 342.29004, 334.9179, 327.46625, 320.25214, 312.79993, 305.1889, 297.5776, 289.966, 282.27484, 274.82126, 267.28812, 259.9926, 252.61752, 245.5594, 238.50105, 231.60107, 224.62155, 217.64178, 210.34451, 203.36426, 196.30444, 189.2444, 182.26343, 175.2029, 168.22147, 161.23978, 154.25786, 147.11702, 140.45201, 133.86613, 127.04199, 120.69374, 114.42466, 107.917305, 101.72719, 95.61626, 89.74323, 83.94942, 78.39354, 72.67877, 67.162285, 61.76471, 56.366997, 51.286663, 45.88867, 39.93484, 34.695328, 29.296898, 24.215893, 19.29355, 13.81532, 8.575136, 3.255418, NaN, NaN, 499.4999, 494.90576, 488.9649, 480.9643, 473.35947, 465.27902, 456.80212, 448.48337, 440.16425, 431.6863, 423.1288, 414.57095, 406.09198, 397.4542, 388.73676, 380.0982, 371.69708, 363.37488, 354.97305, 346.88797, 338.84222, 331.07358, 323.30466, 315.53546, 308.08307, 300.63043, 293.2568, 285.8829, 278.66736, 271.4515, 264.31476, 257.1777, 250.11975, 242.82362, 235.44792, 227.43744, 219.66461, 212.12944, 204.83195, 197.53423, 190.27588, 183.05696, 176.07578, 169.01501, 161.95401, 154.7341, 147.43457, 140.37283, 132.99345, 125.45509, 118.55131, 111.88536, 105.06048, 98.55282, 92.20368, 86.17182, 80.219154, 74.10757, 68.15455, 62.439487, 56.883026, 51.802704, 46.642868, 41.32413, 35.767097, 30.765638, 25.764055, 20.682959, 15.839919, 10.996766, 6.4710927, 2.6599216, NaN, NaN, 498.86676, 493.95575, 487.4604, 478.66754, 469.55743, 460.6846, 451.96985, 443.33392, 434.77692, 426.29877, 418.37494, 410.6093, 402.9226, 395.1564, 386.99362, 379.0683, 371.22192, 363.53378, 355.68683, 347.91882, 340.42798, 333.2143, 326.0004, 318.70694, 311.57178, 304.67426, 297.6179, 290.48203, 283.2666, 276.13022, 268.7557, 261.38095, 254.08519, 246.7892, 239.33432, 231.95848, 224.50307, 217.20602, 210.14668, 202.92844, 195.90826, 189.08617, 182.18451, 175.36195, 168.53918, 161.87485, 155.2103, 148.54555, 141.95992, 135.37407, 128.86736, 122.04304, 115.29784, 108.63178, 102.36231, 96.17201, 90.45773, 84.66392, 78.79057, 72.837685, 67.04337, 61.328274, 55.851154, 50.215126, 44.578945, 39.339535, 34.496933, 29.812996, 25.208344, 20.524193, 16.23691, 12.187729, 7.265085, 3.2951252, NaN, NaN, 499.61975, 494.788, 488.45105, 480.13354, 471.97412, 464.05203, 455.892, 447.89008, 439.80862, 432.04376, 424.35788, 416.59247, 408.7475, 400.90225, 392.8982, 384.9731, 377.0477, 369.35974, 361.35446, 353.58667, 345.77896, 337.9313, 330.16263, 322.2351, 314.30728, 306.617, 298.92642, 291.31485, 283.9409, 276.40805, 268.95422, 261.42087, 253.56999, 245.71883, 237.78804, 230.01558, 222.24283, 214.70773, 207.01373, 199.39876, 192.18013, 184.88193, 177.58347, 170.60208, 163.62045, 156.55927, 149.73584, 142.75351, 135.5329, 128.8675, 122.36057, 115.853455, 109.26676, 102.759224, 96.09275, 89.90226, 83.79095, 77.8382, 71.96465, 66.17031, 60.53456, 54.581135, 49.02445, 43.62638, 37.91062, 32.988594, 28.066444, 23.144178, 17.98361, 13.140498, 8.138474, 3.2951286, NaN, NaN, 500.88742, 496.2933, 490.27325, 481.32208, 472.13287, 462.94324, 454.22855, 445.8304, 437.11502, 428.24078, 419.60385, 411.28357, 402.88367, 394.64197, 386.3999, 377.999, 369.59778, 361.3547, 353.26984, 345.1847, 337.09918, 329.01337, 321.08582, 313.3165, 305.78473, 298.01483, 290.24466, 282.55347, 274.62408, 266.9323, 258.84375, 251.07208, 242.9829, 234.89339, 226.88287, 219.18932, 211.41615, 203.80133, 196.26556, 188.9675, 181.66917, 174.44992, 167.23041, 160.16933, 153.10802, 146.44318, 139.85745, 133.0335, 126.28864, 119.940346, 113.59186, 107.32253, 100.814926, 93.910286, 87.00542, 79.78284, 73.03624, 66.60692, 60.49491, 54.54148, 48.865715, 43.1501, 37.751873, 32.43289, 27.272556, 21.953304, 16.554518, 10.917398, 5.359523, 1.7865233, NaN, NaN, 503.1451, 498.63025, 492.8479, 484.8474, 477.16348, 469.2416, 460.9233, 452.76312, 444.28568, 436.12485, 427.88443, 419.72293, 411.64038, 403.31973, 395.39502, 387.54926, 379.22766, 371.06424, 362.82123, 354.5779, 346.4135, 338.09024, 329.68738, 321.2049, 312.24637, 303.60458, 295.12103, 286.55783, 277.75638, 269.27176, 261.18326, 253.09447, 245.4812, 237.62971, 229.85724, 222.56036, 214.86664, 207.33127, 199.87494, 192.25969, 184.60449, 176.67134, 168.89656, 161.04214, 153.5048, 146.04652, 138.74667, 131.60526, 124.542946, 117.40104, 110.73503, 104.14817, 97.481735, 91.132545, 84.46568, 77.95735, 71.13132, 64.86069, 58.90738, 53.19204, 47.476543, 41.760887, 36.203846, 31.043602, 25.56566, 19.928787, 14.212361, 9.13096, 4.3670316, 1.5880224, NaN, NaN, 499.8978, 495.066, 488.64987, 480.33234, 472.0145, 463.22095, 454.5855, 445.79123, 436.99658, 428.2808, 419.4854, 411.1651, 403.08218, 395.2367, 387.31168, 379.54483, 371.69846, 364.0103, 356.32187, 348.7124, 341.06302, 333.453, 326.1598, 318.86633, 311.5726, 303.9615, 296.66724, 289.21417, 281.7608, 274.54507, 267.01187, 259.47842, 252.02397, 244.72789, 237.35222, 230.13492, 222.75874, 215.30298, 208.00558, 200.6286, 193.29102, 185.91351, 178.53574, 171.1577, 163.7794, 156.55951, 149.65674, 142.99179, 136.16791, 129.66121, 123.15431, 116.72656, 110.37797, 103.949814, 97.759544, 91.8072, 85.61656, 80.21945, 74.74282, 69.26605, 63.947884, 58.629578, 53.311134, 47.59564, 41.72121, 36.32294, 31.242088, 25.922934, 21.31818, 16.95151, 11.790776, 6.788712, 2.977533, NaN, NaN, 503.34363, 498.98718, 493.28406, 484.9667, 476.41138, 467.8557, 459.53732, 450.90173, 442.34497, 433.62943, 424.5173, 415.95944, 407.32202, 398.44647, 389.9668, 381.56604, 373.00644, 364.60498, 356.28244, 348.1181, 339.79492, 331.78845, 323.7817, 315.77466, 307.84656, 299.83887, 292.06873, 284.13974, 276.4483, 268.598, 260.74738, 253.05507, 245.36249, 237.6696, 229.89713, 222.20366, 214.50992, 206.41927, 198.72493, 190.87166, 183.01807, 175.32286, 167.9447, 160.56628, 153.34627, 146.04668, 138.9055, 132.00214, 125.3366, 118.750206, 112.24295, 105.497406, 98.91037, 92.56122, 86.44998, 80.65604, 74.86192, 69.147026, 63.43197, 57.716755, 52.16014, 46.92091, 41.443386, 36.52143, 31.996304, 27.153513, 22.151821, 17.070612, 12.783242, 8.416387, 3.9700367, NaN, NaN, 499.89847, 495.1459, 489.1258, 480.8875, 472.49042, 464.09302, 455.7745, 447.13873, 438.42334, 429.8661, 421.62543, 413.38443, 405.1431, 397.05994, 389.05573, 381.05118, 372.96707, 364.72415, 356.7979, 349.26773, 341.3409, 333.33453, 325.4071, 317.24155, 309.23422, 301.30588, 293.2979, 285.36896, 277.51898, 269.6687, 261.73883, 253.65004, 245.64024, 237.63013, 229.46107, 221.52965, 213.67723, 205.66586, 197.89217, 189.95953, 182.06624, 174.52965, 167.31013, 160.24904, 153.10837, 145.88809, 138.58821, 131.68483, 124.54317, 117.401245, 110.49715, 103.91027, 97.4819, 91.05334, 85.021416, 79.06868, 73.115776, 67.400826, 61.368206, 56.208588, 50.69162, 45.452347, 40.60987, 35.846664, 30.686403, 25.764185, 20.444881, 14.966647, 9.250073, 3.9303396, 1.2307205, NaN, NaN, 500.6909, 496.25516, 490.31433, 482.15527, 474.31277, 466.1531, 457.83466, 449.75357, 441.75137, 433.90735, 425.9838, 418.05994, 410.215, 402.29053, 394.2865, 386.36142, 378.59454, 370.90662, 363.0599, 354.9751, 346.96924, 339.3594, 331.7493, 323.98038, 316.52826, 308.67944, 301.1475, 293.61526, 286.16208, 278.7086, 271.01694, 263.4043, 255.8707, 248.3368, 241.04057, 233.42683, 225.89212, 218.27782, 210.5046, 202.73108, 194.87793, 186.78651, 178.7741, 170.92004, 163.14502, 155.29037, 147.67345, 140.21494, 132.91486, 125.85258, 119.107475, 112.67958, 105.85468, 99.42638, 93.07723, 86.80726, 80.457726, 74.02862, 67.519936, 60.85229, 54.3035, 48.27049, 42.71361, 37.632904, 32.631462, 27.78868, 23.104567, 17.46761, 12.386277, 7.463616, 2.6996372, NaN, NaN, 500.17624, 495.5821, 489.4828, 480.84842, 471.73837, 462.9448, 454.38855, 445.91116, 437.67114, 429.7477, 421.82397, 414.13766, 406.37186, 398.84344, 391.07706, 383.46884, 375.86038, 368.0931, 360.48404, 352.55768, 344.78952, 337.10034, 329.09378, 321.08688, 313.39682, 305.78577, 298.01584, 290.32492, 282.5544, 274.62503, 267.1711, 259.63763, 251.78668, 244.17334, 236.16315, 228.23198, 220.22118, 212.28938, 204.4366, 196.42488, 188.65082, 181.1938, 173.89517, 166.99297, 160.24922, 153.50525, 147.07843, 140.57205, 134.30354, 128.03482, 121.448494, 115.17939, 108.91009, 102.32315, 95.89473, 89.54547, 83.592865, 77.481346, 71.29027, 65.099, 58.7091, 52.596832, 46.643154, 41.006844, 36.08487, 31.87728, 28.145948, 23.144272, 17.824894, 13.537534, 9.329481, 5.438941, 2.104133, NaN, NaN, 499.5824, 494.8298, 488.49286, 480.01685, 471.9366, 464.09372, 455.93365, 447.77322, 439.29556, 430.81757, 422.3392, 413.78125, 405.22296, 396.42657, 387.6298, 378.99115, 370.4314, 361.87128, 353.46936, 345.14636, 336.62485, 327.98407, 319.58075, 311.49423, 303.56595, 295.55807, 287.39133, 279.3828, 271.5326, 263.68207, 255.91057, 248.21806, 240.7632, 233.14944, 225.69403, 218.15903, 210.70308, 203.24684, 195.949, 188.80956, 181.47153, 174.25224, 167.03271, 159.81291, 152.59286, 145.37257, 138.15201, 131.01056, 123.472084, 116.09204, 108.7911, 101.80734, 94.58525, 87.442276, 80.775276, 74.743034, 68.710625, 62.99554, 57.359676, 51.72366, 45.690567, 40.05423, 35.05284, 30.13072, 25.446657, 20.921274, 16.792767, 11.632016, 5.5183425, 1.945332, NaN, NaN, 499.85992, 494.9489, 488.69116, 480.13596, 471.73886, 463.42062, 454.62668, 445.8324, 436.80002, 428.16342, 419.8434, 411.5231, 403.28168, 395.03995, 386.79785, 378.3177, 370.1542, 361.9904, 353.58847, 345.58255, 337.53665, 329.68866, 321.76108, 313.8332, 305.905, 298.0558, 289.9684, 282.35648, 274.74426, 267.13174, 259.67755, 252.22311, 244.927, 237.63063, 230.01675, 222.64053, 215.50201, 208.12527, 200.90692, 193.68832, 186.3108, 178.93301, 171.3963, 163.77997, 156.00467, 148.22906, 140.61188, 133.3118, 126.09081, 118.94893, 111.965515, 105.21995, 98.87097, 92.998, 87.36296, 81.64839, 75.854294, 69.66316, 63.47184, 57.121574, 50.92987, 44.737984, 38.70468, 32.829983, 27.352068, 21.953402, 16.71338, 11.632023, 7.503326, 2.7393415, NaN, NaN, 498.2365, 493.32544, 487.06766, 478.82925, 470.66974, 462.5099, 454.19128, 446.18924, 438.02844, 429.6296, 421.38892, 413.3856, 405.46124, 397.69507, 389.77008, 382.16183, 374.31552, 366.4689, 358.8598, 351.2504, 343.56143, 336.03076, 328.4205, 320.7307, 313.1199, 305.50882, 297.81815, 290.2858, 282.67386, 274.98233, 267.05264, 259.28125, 251.66817, 244.29272, 236.917, 229.54105, 222.24413, 215.10558, 207.96678, 200.90707, 193.72812, 186.50926, 179.05215, 171.6741, 164.21645, 156.75851, 149.6177, 142.87337, 136.20816, 129.62209, 123.27386, 117.08415, 110.57682, 104.62482, 98.59328, 92.561554, 86.609024, 80.65633, 74.8622, 68.82977, 63.233757, 57.677273, 51.961872, 46.643234, 42.277084, 38.149002, 33.94145, 29.654419, 25.3673, 20.68312, 17.030975, 12.267209, 7.900326, 3.2951477, NaN, NaN, 500.53387, 495.9397, 489.84042, 481.91898, 474.2349, 466.15442, 457.83594, 449.75482, 441.67337, 433.5916, 425.27185, 417.42715, 409.50296, 401.7369, 394.1291, 386.20398, 378.27856, 370.35284, 362.34756, 354.0249, 345.66226, 337.49747, 328.936, 320.69125, 312.60477, 304.59723, 296.5101, 288.89838, 281.2071, 273.35693, 265.90298, 258.52805, 251.23215, 243.77737, 236.40164, 229.10497, 221.88733, 214.35219, 206.89607, 199.51901, 191.98305, 184.60545, 177.4656, 170.40483, 163.42316, 156.67928, 149.85582, 143.03215, 136.12889, 128.82864, 121.686844, 114.46545, 107.32315, 100.339325, 93.514, 86.84718, 80.41826, 73.671646, 67.24231, 61.130283, 55.45467, 49.739204, 44.579277, 39.895535, 34.89413, 29.336876, 23.779469, 18.460094, 13.934548, 8.614918, 2.9775472, NaN, NaN, 499.54398, 494.79138, 488.61282, 480.29526, 471.89813, 463.81757, 455.41977, 447.18008, 439.09854, 430.93744, 422.9345, 414.53503, 406.13525, 397.97284, 389.96863, 381.8056, 373.88, 366.11264, 358.18643, 350.3392, 342.4124, 334.24747, 326.08224, 317.99594, 309.98862, 301.981, 293.81445, 285.80618, 277.55972, 269.075, 260.9072, 252.81834, 244.64986, 236.48106, 228.1533, 220.3011, 212.84521, 205.30972, 198.01193, 190.71388, 183.45525, 176.63268, 169.73056, 162.82819, 155.84627, 149.18147, 142.51645, 135.77188, 129.02708, 122.044, 115.21939, 108.79135, 102.680565, 96.887054, 90.93465, 84.823326, 78.71182, 72.67951, 66.56764, 60.931866, 55.653145, 50.3346, 45.492218, 40.729107, 36.204052, 31.758286, 25.407022, 19.690718, 16.117945, 13.497873, 9.289808, 3.414252, NaN, NaN, 498.87097, 494.03912, 487.70212, 479.54297, 471.46268, 463.1444, 454.8258, 446.50687, 438.26685, 430.18494, 422.18198, 414.09943, 406.17508, 398.0127, 389.9292, 381.92468, 374.07834, 365.99393, 358.147, 350.06195, 342.37296, 334.76294, 326.99408, 319.22495, 311.4555, 303.68576, 295.91574, 288.54187, 280.92984, 273.63474, 266.26007, 258.96445, 251.82718, 244.61034, 237.55186, 230.41385, 223.11694, 215.66115, 208.28441, 200.9074, 194.00607, 187.18385, 180.52008, 173.85608, 166.95386, 159.97206, 152.91069, 146.0871, 139.1046, 131.96315, 125.13887, 118.393715, 111.648346, 104.98211, 98.71248, 92.60139, 86.49011, 80.378654, 74.505135, 68.63145, 63.194168, 57.637672, 51.922264, 46.60362, 41.364216, 36.20407, 30.488064, 24.930683, 20.087698, 14.84762, 8.654626, 3.176052, NaN, NaN, 499.9803, 495.3861, 489.44522, 481.6822, 474.0773, 466.15524, 458.3121, 450.231, 441.91187, 433.51315, 425.2726, 416.95245, 408.55276, 400.23193, 391.99005, 383.51007, 375.26752, 366.8661, 358.62286, 350.69638, 342.5714, 334.6443, 326.79614, 318.94772, 311.09897, 303.4878, 295.4799, 287.70953, 279.85962, 272.0094, 264.00027, 255.91151, 247.90176, 240.05031, 232.11925, 224.34651, 216.49417, 208.64151, 200.5506, 192.93532, 185.35942, 177.82292, 170.36546, 162.90775, 155.29108, 147.83281, 140.69167, 133.78831, 126.80539, 119.90157, 112.75945, 105.934525, 99.42683, 92.99829, 86.72829, 80.77557, 75.06081, 69.187126, 63.313286, 57.59803, 51.961998, 46.32581, 41.0864, 35.926243, 31.004124, 25.605536, 20.603777, 15.522498, 10.679288, 5.9947615, 2.580548, NaN, NaN, 499.22815, 494.63397, 488.69302, 481.0884, 473.64194, 466.03674, 458.27283, 450.35016, 442.5064, 434.7416, 427.05576, 419.21112, 411.36618, 403.60022, 395.83395, 387.90887, 380.06277, 372.2956, 364.44888, 356.91895, 349.19055, 341.26367, 333.4158, 325.4883, 317.48126, 309.4739, 301.54553, 293.61682, 285.9257, 278.23428, 270.54257, 263.0092, 255.31693, 247.86229, 240.48668, 233.19012, 226.13126, 219.07214, 211.77483, 204.71523, 197.65538, 190.27797, 182.97963, 175.68103, 168.38217, 161.1624, 154.02171, 146.80142, 139.34285, 131.80464, 124.10746, 116.72741, 109.90261, 103.315674, 97.04598, 90.93483, 85.140976, 79.42632, 73.39402, 67.282166, 61.170124, 55.296047, 49.104267, 43.38861, 37.831573, 33.385834, 30.130854, 26.399473, 21.953485, 17.5074, 12.584836, 7.265157, 2.659951, NaN, NaN, 500.6938, 495.62436, 489.68347, 481.2075, 472.41428, 463.6207, 454.58905, 445.71548, 436.68307, 427.9672, 419.3302, 410.93057, 402.3721, 394.05103, 385.9674, 377.7249, 369.24432, 361.0012, 352.59918, 344.11758, 335.71487, 327.31183, 318.98773, 310.90115, 302.89352, 294.72702, 286.71875, 278.7895, 270.9392, 263.08862, 255.15845, 247.30727, 239.37648, 231.604, 223.6726, 215.82022, 207.88821, 200.27321, 192.65791, 184.963, 177.5058, 169.81032, 162.27324, 154.89456, 147.6743, 140.61249, 133.23303, 126.01201, 119.26688, 112.442154, 105.45849, 98.71268, 92.125374, 85.537865, 79.267624, 73.15594, 67.20283, 61.249535, 55.137314, 49.104294, 43.30925, 37.91098, 32.671345, 27.987318, 23.700148, 19.730465, 16.23708, 11.790869, 6.6299663, 2.8981552, NaN, NaN, 499.82272, 495.14932, 488.97076, 481.2869, 473.7612, 466.23526, 458.62976, 450.78635, 442.78415, 434.94012, 426.85806, 418.7757, 410.61377, 402.2138, 393.73422, 385.41278, 377.09103, 368.6104, 360.36725, 352.12375, 343.9988, 335.75467, 327.5102, 319.1068, 311.0995, 303.0919, 295.24252, 287.39285, 279.6222, 272.08914, 264.4765, 257.0222, 249.40898, 241.79552, 234.41968, 227.0436, 219.66724, 212.44925, 205.38966, 198.2505, 191.26976, 184.20944, 177.22821, 169.9294, 162.63034, 155.41035, 148.26945, 141.20766, 134.14561, 127.24204, 120.10017, 113.11675, 106.529915, 100.65713, 94.70481, 88.83169, 82.9584, 76.926186, 70.97318, 64.94062, 58.78882, 52.835285, 46.881577, 42.197872, 37.831608, 34.020977, 29.892712, 25.526186, 20.36563, 15.20494, 9.964723, 4.8831716, 1.8659412, NaN, NaN, 498.15964, 493.24857, 486.91153, 478.59384, 470.75116, 462.82898, 454.90646, 447.22134, 439.37747, 431.5333, 423.53033, 415.28937, 407.20654, 399.1234, 390.9607, 383.03543, 374.6343, 366.5499, 358.3859, 350.45938, 342.5722, 334.64508, 326.63837, 318.7899, 311.25827, 303.80563, 296.19415, 288.89957, 281.68402, 274.30963, 267.01425, 259.87723, 252.18483, 244.73007, 237.43365, 229.97835, 222.68141, 215.54285, 208.24539, 200.94768, 193.80836, 186.58948, 179.60832, 172.7856, 165.64531, 158.74278, 151.7607, 144.8577, 137.71643, 130.73361, 123.750565, 116.76728, 110.10119, 103.752335, 97.64137, 91.53023, 85.26016, 79.14865, 73.354454, 67.56009, 62.083076, 56.685295, 51.525517, 46.048073, 40.88803, 35.96602, 31.043892, 26.121645, 21.040491, 16.356192, 11.830581, 6.9078717, 2.937859, NaN, NaN, 499.30865, 494.71445, 488.6943, 480.69357, 472.85095, 464.61194, 456.3726, 448.1329, 439.6552, 431.17715, 422.93646, 414.45773, 406.29562, 398.05392, 389.97043, 382.12436, 374.19876, 366.3521, 358.66367, 350.97495, 343.5634, 336.11194, 328.58093, 321.28748, 313.8352, 306.54123, 299.247, 291.71466, 284.49918, 277.12488, 269.7503, 262.61337, 255.39688, 248.33876, 241.43901, 234.53903, 227.16293, 220.10384, 212.88586, 205.66763, 198.21117, 190.91309, 183.53543, 176.3955, 169.41399, 162.5116, 155.45027, 148.3887, 141.72365, 135.13771, 128.55156, 122.04456, 115.61671, 109.1093, 102.83977, 96.411316, 90.141396, 83.79191, 77.75972, 71.96548, 66.29013, 60.81308, 55.41526, 50.176064, 44.85735, 39.856045, 34.854614, 29.932455, 24.930784, 20.008387, 15.324059, 10.401429, 5.558081, 2.0644479, NaN, NaN, 498.87338, 493.88312, 487.54608, 479.06998, 470.11823, 461.16608, 452.1343, 443.3398, 434.70346, 425.98746, 417.35037, 408.8714, 400.70905, 392.3879, 384.14566, 376.06158, 367.97723, 360.1303, 352.20386, 344.1978, 336.11218, 328.02625, 319.78143, 311.69485, 303.92508, 295.7586, 287.82965, 279.9004, 272.05014, 264.51678, 256.58664, 249.0527, 241.4392, 233.7461, 226.29065, 218.6763, 210.90302, 203.36742, 196.22816, 189.24733, 182.4646, 175.95929, 169.53313, 163.10677, 156.83887, 150.25342, 143.66776, 136.84383, 129.86098, 122.71917, 115.73584, 108.672905, 102.0859, 95.65742, 89.62557, 83.355446, 77.56135, 71.84647, 65.97268, 59.93996, 54.224586, 48.11214, 42.15828, 36.759964, 31.758455, 26.836218, 21.993256, 17.229574, 12.465782, 7.3048816, 2.937864, NaN, NaN, 501.4479, 497.01218, 490.99207, 482.99142, 475.54498, 467.62292, 459.93826, 452.09488, 444.40964, 436.4864, 428.56287, 420.55978, 412.79413, 404.9489, 397.3412, 389.57465, 381.72855, 374.04068, 366.2733, 358.50558, 350.89612, 342.89, 335.12143, 327.35254, 319.66266, 313.32025, 307.37408, 301.50702, 295.79837, 290.01025, 284.38058, 278.75076, 273.12076, 267.17343, 261.54312, 255.83336, 250.12344, 244.33405, 238.06863, 231.88235, 225.53725, 219.35059, 213.16373, 206.73872, 200.47217, 194.1261, 187.85915, 181.43335, 174.69002, 167.70845, 160.88531, 154.22064, 147.87314, 141.44609, 135.01884, 128.82945, 122.63987, 116.76753, 110.97438, 104.863625, 98.713, 92.601875, 86.728676, 80.77593, 75.06114, 69.18744, 63.15481, 57.122005, 51.406555, 45.849712, 40.76904, 35.767624, 30.924873, 26.002613, 21.159628, 16.554718, 11.552713, 6.074188, 2.262954, NaN, NaN, 500.93332, 496.41833, 490.47745, 482.2391, 473.68356, 465.28613, 457.20523, 449.12405, 440.9633, 432.9607, 425.03702, 417.1923, 409.34723, 401.73965, 393.73553, 385.81033, 377.8056, 369.80054, 362.1915, 354.89923, 347.3689, 339.8383, 332.06958, 324.45914, 316.76913, 309.07883, 301.46753, 293.61807, 286.00623, 278.23547, 270.46445, 262.53452, 254.6836, 246.91167, 239.13945, 231.129, 223.19756, 215.1865, 207.25443, 199.71869, 192.06367, 184.36871, 176.91147, 169.29527, 162.0755, 154.85547, 147.79388, 140.6527, 133.51126, 126.44893, 119.307, 112.48226, 105.97474, 99.46701, 92.959076, 86.37156, 79.94258, 73.275276, 66.84589, 60.971943, 55.17721, 49.699852, 44.222343, 39.06224, 34.140175, 29.29738, 24.295685, 19.293867, 14.291928, 8.813474, 3.8112786, NaN, NaN, 499.27036, 494.35928, 487.86383, 478.51633, 469.32687, 460.137, 451.34283, 443.18216, 434.54578, 426.22595, 417.6681, 409.42685, 401.50226, 393.65662, 385.9692, 378.28146, 370.51422, 362.82593, 355.13733, 347.607, 339.99713, 332.38696, 324.61798, 317.2451, 309.79263, 302.33994, 295.28342, 287.98877, 280.85245, 273.55728, 266.18256, 258.9662, 251.74956, 244.45335, 237.1569, 230.01883, 222.80118, 215.50395, 208.2858, 201.14671, 194.04704, 187.14545, 180.24362, 173.26224, 166.43929, 160.0128, 153.58612, 147.23859, 141.20825, 135.01904, 128.59157, 122.08456, 115.49798, 109.30798, 103.35589, 97.562355, 92.00676, 86.2129, 80.33951, 74.54532, 68.51284, 62.638943, 56.685497, 51.20817, 46.127625, 41.523266, 36.998196, 32.314243, 27.630186, 22.787233, 17.467793, 11.989418, 6.0344973, 2.2232563, NaN, NaN, 499.19165, 493.7261, 487.46826, 478.59604, 470.11957, 461.5635, 453.24478, 445.00494, 436.52707, 428.44504, 420.20422, 411.88382, 403.7216, 395.55902, 387.55466, 379.4707, 371.4657, 363.4604, 355.45477, 347.7659, 340.0371, 332.50623, 324.89578, 317.68146, 310.3083, 302.7763, 295.24408, 287.47366, 279.54437, 271.6941, 263.84348, 255.91328, 247.98279, 240.21059, 232.59673, 225.22054, 217.76476, 210.38803, 203.40765, 196.34772, 189.60486, 182.78244, 176.03912, 169.21626, 162.31383, 155.64919, 149.14302, 142.47795, 135.97137, 129.22653, 122.48146, 116.21231, 110.339775, 104.30834, 98.43546, 92.562416, 86.6892, 80.73644, 74.70415, 68.59229, 62.361183, 56.566483, 50.851, 45.373516, 40.13404, 35.132603, 30.369213, 25.526321, 20.762707, 15.840191, 10.7587595, 5.7566023, 2.4217627, NaN, NaN, 502.04346, 497.68692, 491.98367, 484.22067, 476.69504, 468.85226, 460.8507, 452.6904, 444.45056, 436.05188, 428.04907, 420.12518, 412.3595, 404.51425, 396.748, 388.98138, 381.69006, 374.16068, 366.78955, 359.25964, 351.61053, 343.92154, 335.99442, 328.22556, 320.21854, 312.29053, 304.60004, 296.7507, 288.82175, 281.2097, 273.51804, 265.74683, 258.0546, 250.44139, 242.90723, 235.6107, 228.55186, 221.41348, 214.03688, 206.58069, 199.48119, 192.42111, 185.59879, 178.85558, 172.03279, 165.05112, 158.0692, 151.08704, 143.62857, 136.48721, 129.74239, 122.75926, 115.45847, 108.55423, 102.04656, 96.014885, 90.14177, 84.34785, 78.791885, 73.23576, 68.116066, 62.877174, 57.161865, 51.20825, 45.25446, 39.3005, 33.981476, 28.900494, 23.898777, 19.055729, 13.974375, 8.416499, 3.414282, NaN, NaN, 499.35052, 494.7563, 488.81534, 481.21063, 473.92255, 466.47577, 458.79105, 451.3437, 443.81686, 436.52747, 429.15857, 421.7894, 414.34073, 407.0503, 399.83884, 392.46863, 385.0189, 377.33112, 369.5638, 361.9547, 354.50388, 346.9735, 339.36362, 331.67413, 324.46002, 317.08713, 309.79324, 302.3405, 295.1254, 287.91, 280.93228, 274.03357, 266.97607, 260.2355, 253.41544, 246.67444, 239.61598, 232.6366, 225.73628, 218.83574, 211.89531, 204.75633, 197.77577, 190.79495, 183.81392, 177.2293, 170.64447, 164.13878, 158.02959, 152.07889, 146.20738, 140.65309, 134.93994, 129.22664, 123.43382, 117.1647, 111.13347, 105.10206, 99.14983, 92.87997, 86.6496, 80.45872, 74.4264, 68.71141, 62.91689, 57.042816, 51.724255, 46.32617, 41.166107, 36.0853, 31.004366, 26.161484, 21.318487, 15.919601, 10.282378, 5.0420027, 1.7071488, NaN, NaN, 500.5391, 496.18253, 490.40002, 482.95383, 475.26968, 467.82294, 460.37595, 452.69098, 445.0057, 437.63712, 430.189, 422.58215, 414.81653, 407.28836, 399.44293, 391.83493, 383.90967, 376.3011, 368.85077, 361.32092, 353.9097, 346.3793, 339.32425, 331.95187, 324.7378, 317.36487, 309.9917, 302.45972, 295.40317, 288.34637, 281.36862, 274.54926, 267.80893, 260.9098, 253.85182, 246.87291, 239.73515, 232.4385, 224.82436, 217.13058, 209.2779, 201.50423, 193.73027, 186.35266, 179.05412, 171.99333, 164.85297, 157.55367, 150.73018, 143.74776, 136.60641, 129.54416, 122.481674, 115.65701, 108.75276, 101.84828, 95.26103, 88.75294, 82.24464, 76.450485, 70.77524, 65.13952, 59.265507, 53.47071, 47.834515, 42.595097, 37.593708, 32.592197, 27.431782, 22.35063, 17.428143, 12.584935, 7.662214, 3.3745856, NaN, NaN, 499.0346, 494.36115, 488.34094, 480.4986, 472.8936, 465.12985, 457.04892, 449.12613, 441.20303, 433.2004, 425.039, 417.1942, 408.9529, 400.86978, 392.8656, 384.94034, 376.69775, 368.61337, 360.52866, 352.83997, 344.75464, 336.8275, 329.13794, 321.3688, 313.67865, 305.9882, 298.45602, 290.9236, 283.70807, 276.2544, 268.80045, 261.2669, 253.81242, 246.5956, 239.45781, 232.16115, 225.1815, 218.51888, 211.38013, 204.08247, 196.78456, 189.48639, 181.94995, 174.73059, 167.43164, 160.52911, 153.309, 145.85059, 138.47125, 131.56776, 124.82276, 118.47431, 112.36375, 106.57044, 100.93571, 95.61827, 90.0626, 84.42741, 78.55394, 72.60094, 66.52869, 60.416573, 54.780563, 49.22378, 44.46071, 39.856297, 35.331173, 30.805946, 26.042444, 21.199434, 16.435709, 11.8306675, 7.0667224, 2.9378805, NaN, NaN, 499.2727, 494.67844, 488.81668, 481.13275, 474.16153, 466.71472, 459.3469, 451.8203, 444.5312, 436.8456, 429.39746, 422.18677, 415.05505, 407.9231, 400.9494, 393.7377, 387.00128, 380.10614, 373.21075, 366.31512, 359.49857, 352.52322, 345.46835, 338.57184, 331.59576, 324.38165, 317.24655, 310.11124, 302.7378, 295.04694, 287.75223, 280.5366, 273.24136, 266.1045, 258.80878, 251.4335, 244.13727, 236.84077, 229.86127, 222.80222, 215.78258, 208.88168, 201.74258, 194.99988, 188.25694, 181.59312, 175.16708, 168.50284, 161.6797, 154.69765, 147.636, 140.81216, 134.46422, 128.11606, 122.16448, 116.45081, 110.578255, 104.705536, 98.91201, 93.277054, 87.641945, 81.68919, 75.974396, 70.25943, 64.70307, 59.384693, 54.54247, 49.858894, 45.095833, 40.332657, 35.01365, 29.376934, 23.263702, 17.229687, 10.877897, 4.9229155, 1.6674525, NaN, NaN, 499.74823, 495.23322, 489.45068, 481.21225, 472.8943, 464.81363, 456.7327, 448.49295, 440.41138, 432.32947, 424.64343, 416.7194, 408.79504, 401.18738, 393.42093, 385.57495, 377.57016, 369.56503, 361.87668, 354.6636, 347.48993, 340.11783, 332.98328, 325.92773, 318.71344, 311.57812, 304.3633, 296.7518, 289.0607, 281.6072, 274.15344, 266.5408, 259.0072, 251.23538, 243.30467, 235.69089, 227.83888, 220.0659, 212.5306, 204.91566, 197.37979, 189.68498, 182.06923, 174.45317, 167.1542, 160.33101, 153.42824, 146.28722, 139.46333, 132.71857, 126.13229, 119.783875, 113.3559, 106.848366, 100.73744, 94.86444, 89.22937, 83.4354, 77.72065, 72.00573, 65.93346, 59.821316, 54.423428, 49.660465, 44.897392, 40.292988, 35.609085, 30.92508, 26.39975, 21.556742, 16.396034, 10.44121, 4.248009, 0.9131309, NaN, NaN, 500.4615, 495.6296, 489.45102, 480.89572, 472.41928, 463.6256, 455.14847, 446.5125, 438.11392, 429.71497, 421.55338, 413.15375, 404.83304, 396.03647, 387.7943, 379.47256, 371.46753, 363.2244, 355.21872, 347.292, 339.00824, 331.0809, 322.83615, 314.82892, 306.97992, 299.44778, 291.5982, 283.82764, 276.05676, 268.52347, 261.06924, 253.77333, 246.15994, 239.18074, 231.96338, 224.58711, 217.28992, 209.7545, 202.2188, 194.52415, 187.14656, 179.61003, 171.99388, 164.61548, 157.55417, 150.33394, 143.11343, 135.97205, 128.8304, 121.76786, 114.62572, 107.80077, 101.05497, 94.54704, 88.11827, 81.76867, 75.49825, 69.22764, 63.194965, 57.71778, 52.359528, 46.80267, 41.24566, 35.76789, 30.686928, 25.526447, 20.28644, 15.125697, 9.726626, 4.3274136, 1.2307415, NaN, NaN, 500.42236, 495.43207, 489.09503, 481.015, 473.41, 465.01248, 456.8523, 449.16718, 441.48175, 434.03375, 426.50626, 419.29544, 412.08438, 404.9523, 397.81998, 390.84592, 383.87164, 376.50082, 369.28824, 361.9962, 354.46603, 347.17343, 339.56348, 332.03253, 324.5013, 317.12836, 309.91373, 302.61954, 295.72156, 288.74402, 281.52838, 274.55038, 267.49286, 260.51437, 253.13914, 246.00156, 238.86374, 231.72566, 224.66666, 217.6074, 209.99266, 202.61562, 195.47629, 188.25737, 181.19687, 174.5328, 167.78918, 161.12468, 154.22194, 147.23961, 140.3364, 133.3536, 126.21186, 119.62537, 113.435455, 107.48344, 101.45189, 95.81699, 89.70573, 83.514915, 77.32391, 71.13272, 65.02073, 58.908546, 52.95495, 47.55687, 42.873127, 38.030502, 33.02898, 27.550985, 22.231632, 17.626707, 12.227696, 6.9873447, 3.0172918, NaN, NaN, 499.59106, 495.07602, 488.9766, 481.3719, 474.2422, 466.71616, 459.18985, 451.66324, 444.13638, 436.53, 428.68564, 420.99945, 413.23373, 405.54697, 398.01843, 390.1726, 382.40573, 374.7178, 366.95035, 359.26187, 351.692, 344.16147, 336.63068, 329.1789, 321.64755, 313.7988, 306.10834, 298.73474, 291.20227, 283.66956, 276.53302, 269.47556, 262.17993, 255.28058, 248.38098, 241.48117, 234.42249, 227.76015, 221.09758, 214.11752, 206.97859, 199.5221, 192.38264, 185.00496, 177.46834, 170.01077, 162.94965, 155.9676, 149.06468, 142.32022, 135.49619, 128.90999, 122.64099, 115.89566, 108.832664, 102.404335, 95.7377, 89.30896, 83.118126, 77.08585, 71.25185, 65.377975, 59.742085, 54.026653, 48.549213, 43.2304, 38.38778, 33.545044, 28.54341, 23.382866, 18.142796, 13.140785, 8.376852, 3.8510122, NaN}
    CHLA = 
      {NaN, 0.168, 0.17700000000000002, 0.195, 0.18, 0.168, 0.17400000000000002, 0.189, 0.171, 0.168, 0.171, 0.30300000000000005, 0.17400000000000002, 0.17400000000000002, 0.17700000000000002, 0.17400000000000002, 0.171, 0.18, 0.183, 0.17400000000000002, 0.165, 0.183, 0.18, 0.183, 0.17400000000000002, 0.18, 0.003, 0.18, 0.183, 0.195, 0.186, 0.17700000000000002, 0.186, 0.186, 0.183, 0.195, 0.186, 0.003, 0.201, 0.21000000000000002, 0.23099999999999998, 0.23399999999999999, 0.261, 0.273, 0.264, 0.28200000000000003, 0.29700000000000004, 0.31200000000000006, 0.318, 0.318, 0.315, 0.321, 0.315, 0.336, 0.327, 0.342, 0.35400000000000004, 0.399, 0.378, 0.375, 0.45899999999999996, 0.513, 0.5880000000000001, 0.678, 0.765, 0.7140000000000001, 0.948, 0.759, 0.795, 0.8130000000000001, 0.921, 0.8400000000000001, 0.927, 0.9450000000000001, 0.8999999999999999, 0.9810000000000001, 0.8640000000000001, 0.9179999999999999, 0.8250000000000001, 0.8160000000000001, NaN, NaN, 0.17400000000000002, 0.17700000000000002, 0.17400000000000002, 0.17400000000000002, 0.17700000000000002, 0.168, 0.171, 0.17400000000000002, 0.171, 0.171, 0.171, 0.168, 0.183, 0.17400000000000002, 0.168, 0.17700000000000002, 0.17700000000000002, 0.171, 0.17700000000000002, 0.17700000000000002, 0.192, 0.17700000000000002, 0.17700000000000002, 0.18, 0.183, 0.17700000000000002, 0.171, 0.17400000000000002, 0.18, 0.20400000000000001, 0.17400000000000002, 0.186, 0.18, 0.18, 0.17700000000000002, 0.195, 0.183, 0.201, 0.17700000000000002, 0.186, 0.186, 0.195, 0.201, 0.22799999999999998, 0.23399999999999999, 0.237, 0.246, 0.249, 0.246, 0.255, 0.273, 0.28200000000000003, 0.30300000000000005, 0.30600000000000005, 0.321, 0.339, 0.327, 0.33, 0.339, 0.39, 0.41700000000000004, 0.579, 0.678, 0.789, 0.75, 0.72, 0.8130000000000001, 0.795, 0.9059999999999999, 0.8640000000000001, 0.867, 0.873, 0.8640000000000001, 0.942, 0.9059999999999999, 0.9359999999999999, 0.9450000000000001, 0.8699999999999999, 0.756, 0.747, 0.72, NaN, NaN, 0.168, 0.168, 0.168, 0.168, 0.168, 0.168, 0.168, 0.168, 0.084, 0.168, 0.171, 0.171, 0.171, 0.171, 0.17700000000000002, 0.171, 0.17700000000000002, 0.17400000000000002, 0.17400000000000002, 0.17400000000000002, 0.18, 0.17400000000000002, 0.17700000000000002, 0.18, 0.17400000000000002, 0.192, 0.186, 0.21600000000000003, 0.243, 0.276, 0.318, 0.366, 0.36, 0.41400000000000003, 0.723, 0.783, 0.909, 0.927, 0.8999999999999999, 0.903, 0.897, 0.9810000000000001, 1.0350000000000001, 1.0290000000000001, 0.942, 0.8370000000000001, 0.687, NaN, NaN, 0.171, 0.171, 0.168, 0.168, 0.168, 0.17400000000000002, 0.165, 0.168, 0.081, 0.18, 0.171, 0.168, 0.168, 0.165, 0.171, 0.168, 0.168, 0.171, 0.168, 0.171, 0.17400000000000002, 0.168, 0.17400000000000002, 0.18, 0.17400000000000002, 0.18, 0.186, 0.18, 0.186, 0.192, 0.21000000000000002, 0.24, 0.252, 0.28200000000000003, 0.324, 0.35400000000000004, 0.192, 0.6120000000000001, 0.66, 0.8280000000000001, 1.0110000000000001, 0.9690000000000001, 1.0410000000000001, 1.131, 1.0410000000000001, 1.0979999999999999, 1.191, 1.059, 0.8550000000000001, 0.645, NaN, NaN, 0.162, 0.165, 0.168, 0.168, 0.165, 0.165, 0.171, 0.162, 0.171, 0.165, 0.165, 0.165, 0.162, 0.168, 0.168, 0.17400000000000002, 0.17400000000000002, 0.168, 0.171, 0.17400000000000002, 0.171, 0.17400000000000002, 0.17700000000000002, 0.168, 0.168, 0.171, 0.18, 0.198, 0.17700000000000002, 0.186, 0.186, 0.20700000000000002, 0.23399999999999999, 0.264, 0.28200000000000003, 0.315, 0.339, 0.41700000000000004, 0.534, 0.687, 0.8220000000000001, 0.474, 1.044, 1.1099999999999999, 0.534, 1.116, 1.158, 1.344, 1.068, 0.786, 0.6000000000000001, 0.51, NaN, NaN, 0.168, 0.162, 0.162, 0.162, 0.165, 0.162, 0.165, 0.165, 0.165, 0.165, 0.165, 0.171, 0.159, 0.165, 0.165, 0.165, 0.165, 0.168, 0.171, 0.165, 0.168, 0.17700000000000002, 0.201, 0.165, 0.168, 0.168, 0.17700000000000002, 0.168, 0.17400000000000002, 0.18, 0.192, 0.192, 0.189, 0.195, 0.195, 0.22799999999999998, 0.132, 0.29700000000000004, 0.33, 0.321, 0.34500000000000003, 0.21300000000000002, 0.507, 0.579, 0.663, 0.9870000000000001, 1.113, 1.305, 1.257, 0.567, 0.891, 0.771, 0.399, 0.639, 0.567, 0.471, NaN, NaN, 0.168, 0.162, 0.162, 0.162, 0.165, 0.162, 0.162, 0.165, 0.162, 0.168, 0.162, 0.165, 0.17400000000000002, 0.165, 0.165, 0.165, 0.162, 0.165, 0.159, 0.162, 0.162, 0.165, 0.168, 0.183, 0.165, 0.168, 0.17400000000000002, 0.168, 0.17700000000000002, 0.17400000000000002, 0.18, 0.183, 0.189, 0.096, 0.198, 0.192, 0.198, 0.22799999999999998, 0.258, 0.29400000000000004, 0.315, 0.324, 0.336, 0.35700000000000004, 0.35400000000000004, 0.43499999999999994, 0.558, 0.687, 1.038, 1.1400000000000001, 1.05, 0.8550000000000001, 0.8460000000000001, 0.735, 0.72, 0.6240000000000001, NaN, NaN, 0.159, 0.159, 0.162, 0.159, 0.168, 0.159, 0.159, 0.162, 0.081, 0.15300000000000002, 0.159, 0.159, 0.162, 0.159, 0.162, 0.159, 0.162, 0.162, 0.165, 0.171, 0.165, 0.171, 0.17400000000000002, 0.165, 0.171, 0.165, 0.17700000000000002, 0.168, 0.17700000000000002, 0.17700000000000002, 0.17400000000000002, 0.195, 0.10800000000000001, 0.23099999999999998, 0.243, 0.258, 0.28800000000000003, 0.29700000000000004, 0.162, 0.339, 0.35100000000000003, 0.339, 0.363, 0.35700000000000004, 0.375, 0.399, 0.405, 0.45299999999999996, 0.45899999999999996, 0.279, 0.753, 0.765, 0.807, 0.405, 0.8130000000000001, 0.747, NaN, NaN, 0.159, 0.159, 0.159, 0.162, 0.15600000000000003, 0.159, 0.162, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.159, 0.159, 0.07800000000000001, 0.165, 0.15600000000000003, 0.159, 0.159, 0.162, 0.162, 0.162, 0.165, 0.159, 0.159, 0.168, 0.162, 0.162, 0.162, 0.168, 0.168, 0.168, 0.165, 0.171, 0.18, 0.195, 0.21600000000000003, 0.23399999999999999, 0.23399999999999999, 0.255, 0.28500000000000003, 0.333, 0.17700000000000002, 0.372, 0.387, 0.375, 0.195, 0.42900000000000005, 0.43499999999999994, 0.44099999999999995, 0.44699999999999995, 0.24, 0.519, 0.522, 0.753, 0.729, 0.789, 0.8340000000000001, 0.777, 0.723, 0.8130000000000001, 0.6990000000000001, NaN, NaN, 0.162, 0.159, 0.15600000000000003, 0.159, 0.159, 0.15600000000000003, 0.15300000000000002, 0.159, 0.084, 0.15600000000000003, 0.159, 0.159, 0.15300000000000002, 0.159, 0.15600000000000003, 0.15600000000000003, 0.159, 0.081, 0.15600000000000003, 0.159, 0.081, 0.162, 0.165, 0.162, 0.15600000000000003, 0.159, 0.162, 0.165, 0.171, 0.171, 0.20700000000000002, 0.17700000000000002, 0.201, 0.22799999999999998, 0.22799999999999998, 0.24, 0.243, 0.246, 0.264, 0.264, 0.258, 0.28200000000000003, 0.29400000000000004, 0.324, 0.34800000000000003, 0.36, 0.381, 0.39, 0.399, 0.393, 0.39, 0.41100000000000003, 0.45899999999999996, 0.675, 0.8370000000000001, 0.78, 0.759, 0.7110000000000001, 0.72, 0.6990000000000001, 0.729, 0.0, NaN, NaN, 0.162, 0.159, 0.15600000000000003, 0.165, 0.15600000000000003, 0.159, 0.159, 0.15300000000000002, 0.081, 0.15600000000000003, 0.162, 0.15600000000000003, 0.159, 0.081, 0.07800000000000001, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.159, 0.162, 0.162, 0.159, 0.165, 0.165, 0.162, 0.165, 0.171, 0.168, 0.168, 0.171, 0.195, 0.21300000000000002, 0.11399999999999999, 0.11699999999999999, 0.21899999999999997, 0.22799999999999998, 0.261, 0.279, 0.279, 0.279, 0.30300000000000005, 0.327, 0.363, 0.393, 0.399, 0.393, 0.41700000000000004, 0.45299999999999996, 0.489, 0.663, 0.6990000000000001, 0.381, 0.795, 0.8130000000000001, 0.8370000000000001, 0.897, 1.008, 0.933, NaN, NaN, 0.159, 0.15300000000000002, 0.162, 0.159, 0.159, 0.15600000000000003, 0.15600000000000003, 0.162, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.081, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.159, 0.15600000000000003, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.165, 0.168, 0.165, 0.168, 0.165, 0.168, 0.168, 0.165, 0.171, 0.168, 0.18, 0.189, 0.21300000000000002, 0.20700000000000002, 0.22199999999999998, 0.21300000000000002, 0.22799999999999998, 0.249, 0.276, 0.321, 0.324, 0.35100000000000003, 0.34500000000000003, 0.198, 0.396, 0.405, 0.41400000000000003, 0.45299999999999996, 0.501, 0.5309999999999999, 0.591, 0.603, 0.66, 0.72, 0.81, 0.8160000000000001, 0.42000000000000004, 0.786, NaN, NaN, 0.159, 0.159, 0.159, 0.159, 0.159, 0.15600000000000003, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.165, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.162, 0.165, 0.17400000000000002, 0.186, 0.201, 0.23099999999999998, 0.22499999999999998, 0.273, 0.34500000000000003, 0.35700000000000004, 0.372, 0.387, 0.43799999999999994, 0.486, 0.5549999999999999, 0.615, 0.759, 0.777, 0.6900000000000001, 0.7110000000000001, NaN, NaN, 0.159, 0.162, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.162, 0.123, 0.165, 0.17400000000000002, 0.17400000000000002, 0.17700000000000002, 0.17700000000000002, 0.186, 0.15300000000000002, 0.21000000000000002, 0.23399999999999999, 0.267, 0.237, 0.375, 0.396, 0.44999999999999996, 0.46199999999999997, 0.519, 0.66, 0.765, 0.729, 0.657, NaN, NaN, 0.159, 0.159, 0.159, 0.15300000000000002, 0.15600000000000003, 0.159, 0.15600000000000003, 0.11699999999999999, 0.162, 0.15600000000000003, 0.15600000000000003, 0.17700000000000002, 0.11699999999999999, 0.11699999999999999, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.159, 0.159, 0.162, 0.12, 0.162, 0.165, 0.126, 0.17400000000000002, 0.17700000000000002, 0.195, 0.201, 0.201, 0.21300000000000002, 0.22199999999999998, 0.237, 0.279, 0.372, 0.324, 0.315, 0.42600000000000005, 0.46199999999999997, 0.483, 0.657, 0.741, 0.642, NaN, NaN, 0.15600000000000003, 0.159, 0.15600000000000003, 0.159, 0.15600000000000003, 0.159, 0.11699999999999999, 0.168, 0.15600000000000003, 0.159, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.159, 0.165, 0.162, 0.165, 0.18, 0.195, 0.21899999999999997, 0.23099999999999998, 0.261, 0.31200000000000006, 0.35400000000000004, 0.405, 0.41400000000000003, 0.405, 0.5369999999999999, 0.639, 0.6930000000000001, 0.6900000000000001, 0.681, 0.519, 0.72, NaN, NaN, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.11399999999999999, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.11699999999999999, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.11699999999999999, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.159, 0.126, 0.171, 0.168, 0.168, 0.171, 0.17400000000000002, 0.189, 0.20400000000000001, 0.21899999999999997, 0.23099999999999998, 0.28200000000000003, 0.30600000000000005, 0.35700000000000004, 0.42300000000000004, 0.41700000000000004, 0.567, 0.6180000000000001, 0.672, 0.729, 0.567, 0.507, NaN, NaN, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15000000000000002, 0.159, 0.162, 0.123, 0.159, 0.162, 0.159, 0.165, 0.165, 0.17400000000000002, 0.138, 0.192, 0.20400000000000001, 0.21899999999999997, 0.22499999999999998, 0.23399999999999999, 0.255, 0.30600000000000005, 0.336, 0.366, 0.42900000000000005, 0.486, 0.5940000000000001, 0.633, 0.678, 0.6960000000000001, 0.759, 0.8370000000000001, 0.6990000000000001, NaN, NaN, 0.15600000000000003, 0.159, 0.159, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.159, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.11399999999999999, 0.11399999999999999, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.12, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.159, 0.162, 0.162, 0.168, 0.165, 0.168, 0.168, 0.171, 0.17700000000000002, 0.138, 0.201, 0.21000000000000002, 0.189, 0.24, 0.261, 0.27, 0.342, 0.43799999999999994, 0.46799999999999997, 0.483, 0.558, 0.513, 0.753, 0.7140000000000001, 0.762, 0.795, 0.8460000000000001, 0.7110000000000001, NaN, NaN, 0.159, 0.15600000000000003, 0.159, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.12, 0.159, 0.15600000000000003, 0.12, 0.162, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.11699999999999999, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.11399999999999999, 0.12, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.11699999999999999, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.159, 0.162, 0.165, 0.171, 0.168, 0.171, 0.183, 0.189, 0.20400000000000001, 0.23399999999999999, 0.23399999999999999, 0.249, 0.273, 0.30000000000000004, 0.366, 0.43499999999999994, 0.507, 0.522, 0.6000000000000001, 0.726, 0.798, 0.723, 0.768, 0.8280000000000001, 0.78, 0.795, 0.636, NaN, NaN, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.11699999999999999, 0.15300000000000002, 0.159, 0.11699999999999999, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.15300000000000002, 0.11399999999999999, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.11399999999999999, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.162, 0.168, 0.171, 0.171, 0.171, 0.17700000000000002, 0.135, 0.186, 0.21000000000000002, 0.22199999999999998, 0.249, 0.252, 0.28500000000000003, 0.327, 0.393, 0.492, 0.552, 0.597, 0.663, 0.51, 0.7080000000000001, 0.7050000000000001, 0.5820000000000001, 0.738, 0.753, 0.657, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.11399999999999999, 0.15600000000000003, 0.15300000000000002, 0.11399999999999999, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.11399999999999999, 0.15300000000000002, 0.11399999999999999, 0.15300000000000002, 0.15300000000000002, 0.159, 0.165, 0.126, 0.171, 0.17400000000000002, 0.18, 0.17700000000000002, 0.186, 0.198, 0.201, 0.22799999999999998, 0.243, 0.264, 0.28200000000000003, 0.339, 0.41400000000000003, 0.36, 0.729, 0.6930000000000001, 0.738, 0.8340000000000001, 0.8340000000000001, 0.7020000000000001, 0.9299999999999999, 0.9179999999999999, 0.768, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11399999999999999, 0.15300000000000002, 0.11399999999999999, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11699999999999999, 0.159, 0.162, 0.129, 0.17700000000000002, 0.186, 0.18, 0.192, 0.198, 0.22199999999999998, 0.22799999999999998, 0.252, 0.30000000000000004, 0.336, 0.42000000000000004, 0.43799999999999994, 0.384, 0.636, 0.738, 0.81, 0.8640000000000001, 0.738, 1.17, 1.158, 0.726, 0.684, NaN, NaN, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.11699999999999999, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.11399999999999999, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.14700000000000002, 0.11399999999999999, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.162, 0.165, 0.165, 0.168, 0.18, 0.249, 0.21000000000000002, 0.22499999999999998, 0.246, 0.264, 0.29400000000000004, 0.33, 0.369, 0.42300000000000004, 0.44399999999999995, 0.501, 0.5700000000000001, 0.6180000000000001, 0.687, 0.8250000000000001, 1.0979999999999999, 1.242, 1.095, 0.8430000000000001, 1.191, NaN, NaN, 0.15600000000000003, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.11399999999999999, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.11399999999999999, 0.11399999999999999, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.123, 0.126, 0.165, 0.171, 0.18, 0.159, 0.22499999999999998, 0.249, 0.261, 0.28500000000000003, 0.35100000000000003, 0.387, 0.387, 0.399, 0.471, 0.519, 0.45899999999999996, 0.8430000000000001, 0.9870000000000001, 0.885, 0.909, 0.903, 0.933, 0.675, 0.9510000000000001, NaN, NaN, 0.15300000000000002, 0.159, 0.15600000000000003, 0.15300000000000002, 0.11699999999999999, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11399999999999999, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.11699999999999999, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.17400000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.11399999999999999, 0.14700000000000002, 0.15000000000000002, 0.11399999999999999, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.11399999999999999, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.168, 0.165, 0.17700000000000002, 0.14100000000000001, 0.20400000000000001, 0.21600000000000003, 0.23099999999999998, 0.237, 0.27, 0.252, 0.36, 0.333, 0.393, 0.5489999999999999, 0.8490000000000001, 0.807, 0.777, 0.789, 0.8640000000000001, 0.8160000000000001, 1.0859999999999999, 1.1400000000000001, 0.9690000000000001, 0.9179999999999999, 0.8610000000000001, 0.9990000000000001, NaN, NaN, 0.159, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.12, 0.15600000000000003, 0.15000000000000002, 0.15000000000000002, 0.11699999999999999, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.11099999999999999, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.11399999999999999, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.162, 0.168, 0.17400000000000002, 0.14100000000000001, 0.192, 0.201, 0.21300000000000002, 0.21300000000000002, 0.21000000000000002, 0.21600000000000003, 0.22499999999999998, 0.24, 0.201, 0.29400000000000004, 0.324, 0.315, 0.363, 0.471, 0.66, 0.732, 0.642, 0.7080000000000001, 1.104, 1.182, 1.104, 1.1099999999999999, NaN, NaN, 0.15300000000000002, 0.159, 0.15600000000000003, 0.15300000000000002, 0.132, 0.15600000000000003, 0.15600000000000003, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.129, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.183, 0.183, 0.189, 0.201, 0.21000000000000002, 0.22499999999999998, 0.237, 0.258, 0.273, 0.28800000000000003, 0.369, 0.43200000000000005, 0.486, 0.5489999999999999, 0.8490000000000001, 0.681, 0.7080000000000001, 0.9059999999999999, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.159, 0.165, 0.183, 0.189, 0.20400000000000001, 0.24, 0.264, 0.276, 0.327, 0.43799999999999994, 0.5880000000000001, 0.789, 0.768, 0.7050000000000001, 0.627, NaN, NaN, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.126, 0.138, 0.17400000000000002, 0.21600000000000003, 0.27, 0.24, 0.318, 0.36, 0.46799999999999997, 0.789, 0.519, 0.759, 0.5820000000000001, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.123, 0.123, 0.126, 0.14700000000000002, 0.123, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.17700000000000002, 0.18, 0.201, 0.261, 0.273, 0.30900000000000005, 0.363, 0.546, 0.615, 0.8280000000000001, 0.8460000000000001, 0.651, 0.507, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.162, 0.198, 0.189, 0.249, 0.276, 0.315, 0.40800000000000003, 0.5820000000000001, 0.5489999999999999, 0.732, 0.603, 0.504, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.123, 0.15600000000000003, 0.183, 0.22799999999999998, 0.249, 0.375, 0.45599999999999996, 0.522, 0.5820000000000001, 0.741, 0.585, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.165, 0.21600000000000003, 0.258, 0.28200000000000003, 0.31200000000000006, 0.387, 0.41700000000000004, 0.723, 0.771, 0.747, 0.8819999999999999, NaN, NaN, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.15300000000000002, 0.159, 0.195, 0.23099999999999998, 0.267, 0.336, 0.48, 0.603, 0.753, 0.909, 0.8340000000000001, 0.6990000000000001, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.126, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.12, 0.14700000000000002, 0.129, 0.17400000000000002, 0.198, 0.246, 0.23399999999999999, 0.321, 0.519, 0.6000000000000001, 0.6960000000000001, 0.909, 0.8999999999999999, 0.8759999999999999, 0.8400000000000001, 0.522, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.126, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.192, 0.237, 0.255, 0.28500000000000003, 0.34800000000000003, 0.654, 0.8939999999999999, 0.978, 0.927, 0.978, 0.738, 0.519, NaN, NaN, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.12, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.162, 0.18, 0.20400000000000001, 0.252, 0.276, 0.24, 0.36, 0.44399999999999995, 0.9239999999999999, 1.092, 1.05, 1.02, 0.942, 0.651, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.15300000000000002, 0.14700000000000002, 0.159, 0.165, 0.171, 0.201, 0.249, 0.273, 0.369, 0.5549999999999999, 1.0470000000000002, 1.071, 0.867, 0.984, 0.7170000000000001, 0.5700000000000001, NaN, NaN, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.15000000000000002, 0.12, 0.162, 0.14400000000000002, 0.20400000000000001, 0.258, 0.30600000000000005, 0.8939999999999999, 1.1219999999999999, 0.8580000000000001, 0.744, 0.8580000000000001, 1.02, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.126, 0.17400000000000002, 0.18, 0.198, 0.22199999999999998, 0.18, 0.23399999999999999, 0.29400000000000004, 0.30000000000000004, 0.378, 0.8819999999999999, 1.1640000000000001, 0.8759999999999999, 0.762, 0.657, 0.723, NaN, NaN, 0.15000000000000002, 0.15600000000000003, 0.15600000000000003, 0.15000000000000002, 0.15600000000000003, 0.15600000000000003, 0.162, 0.18, 0.198, 0.21600000000000003, 0.276, 0.276, 0.9119999999999999, 1.0859999999999999, 0.8340000000000001, 0.768, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.126, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.20700000000000002, 0.18, 0.171, 0.243, 0.30600000000000005, 0.369, 1.143, 1.089, 0.8190000000000001, NaN, NaN, 0.15600000000000003, 0.162, 0.15600000000000003, 0.162, 0.15000000000000002, 0.15000000000000002, 0.132, 0.168, 0.168, 0.186, 0.21000000000000002, 0.23399999999999999, 0.28800000000000003, 0.396, 0.6120000000000001, 1.092, 0.972, NaN, NaN, 0.15600000000000003, 0.162, 0.15000000000000002, 0.15600000000000003, 0.15600000000000003, 0.15000000000000002, 0.15600000000000003, 0.162, 0.168, 0.138, 0.186, 0.198, 0.192, 0.276, 0.46799999999999997, 0.552, 0.972, 0.8340000000000001, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.162, 0.126, 0.15600000000000003, 0.135, 0.168, 0.18, 0.186, 0.22499999999999998, 0.252, 0.29400000000000004, 0.35700000000000004, 0.54, 0.783, 0.663, 1.002, 1.0859999999999999, 0.9299999999999999, 0.6900000000000001, NaN, NaN, 0.165, 0.15300000000000002, 0.159, 0.15300000000000002, 0.135, 0.159, 0.15300000000000002, 0.165, 0.195, 0.30900000000000005, 0.591, 0.777, 0.9870000000000001, 1.0290000000000001, 0.315, NaN, NaN, 0.15600000000000003, 0.159, 0.15300000000000002, 0.15600000000000003, 0.129, 0.15300000000000002, 0.168, 0.20700000000000002, 0.23399999999999999, 0.477, 0.8250000000000001, 0.771, 0.984, 1.059, 0.8280000000000001, NaN, NaN, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.15300000000000002, 0.15300000000000002, 0.165, 0.201, 0.20700000000000002, 0.23099999999999998, 0.43499999999999994, 0.867, 0.903, 1.0470000000000002, 0.879, NaN, NaN, 0.15600000000000003, 0.15000000000000002, 0.126, 0.15600000000000003, 0.162, 0.15600000000000003, 0.15000000000000002, 0.15600000000000003, 0.138, 0.21600000000000003, 0.33, 0.8879999999999999, 0.8939999999999999, 1.002, 0.8939999999999999, NaN, NaN, 0.159, 0.168, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.17400000000000002, 0.17700000000000002, 0.264, 0.5760000000000001, 0.765, 1.0230000000000001, 0.666, 0.477, NaN, NaN, 0.159, 0.159, 0.15300000000000002, 0.162, 0.15300000000000002, 0.15300000000000002, 0.15000000000000002, 0.126, 0.159, 0.186, 0.252, 0.372, 0.591, 0.7170000000000001, 1.008, 0.933, 0.795, NaN, NaN, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.165, 0.21899999999999997, 0.201, 0.31200000000000006, 0.633, 0.8520000000000001, 0.735, NaN, NaN, 0.165, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.129, 0.159, 0.15600000000000003, 0.162, 0.22499999999999998, 0.22799999999999998, 0.264, 0.636, 0.9510000000000001, 0.9630000000000001, 1.026, NaN, NaN, 0.15300000000000002, 0.159, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.21300000000000002, 0.24, 0.366, 0.654, 0.786, 0.933, 0.7140000000000001, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.165, 0.195, 0.21899999999999997, 0.315, 0.44699999999999995, 0.8250000000000001, 0.9390000000000001, 0.933, NaN, NaN, 0.15600000000000003, 0.162, 0.132, 0.15600000000000003, 0.15000000000000002, 0.15000000000000002, 0.132, 0.168, 0.192, 0.21600000000000003, 0.246, 0.384, 0.42000000000000004, 0.8460000000000001, 0.8699999999999999, 1.002, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.159, 0.15300000000000002, 0.132, 0.162, 0.165, 0.21000000000000002, 0.27, 0.42900000000000005, 0.636, 0.765, 0.798, 1.0619999999999998, NaN, NaN, 0.15300000000000002, 0.15600000000000003, 0.129, 0.15300000000000002, 0.132, 0.15600000000000003, 0.165, 0.195, 0.243, 0.28200000000000003, 0.627, 0.6180000000000001, 0.8220000000000001, 1.113, NaN, NaN, 0.15600000000000003, 0.162, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.132, 0.165, 0.189, 0.23099999999999998, 0.24, 0.43799999999999994, 0.621, 0.8550000000000001, 0.9630000000000001, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15300000000000002, 0.135, 0.162, 0.14700000000000002, 0.186, 0.21000000000000002, 0.342, 0.534, 0.8130000000000001, 1.107, 0.774, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.162, 0.162, 0.18, 0.168, 0.22199999999999998, 0.252, 0.402, 0.732, 1.002, 0.504, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.162, 0.168, 0.17400000000000002, 0.21000000000000002, 0.21300000000000002, 0.28200000000000003, 0.45899999999999996, 0.6060000000000001, 0.8400000000000001, 0.51, NaN, NaN, 0.159, 0.159, 0.15300000000000002, 0.159, 0.159, 0.15300000000000002, 0.159, 0.171, 0.21300000000000002, 0.261, 0.35700000000000004, 0.741, 0.9510000000000001, 0.483, NaN, NaN, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.159, 0.159, 0.18, 0.201, 0.31200000000000006, 0.45899999999999996, 0.768, 0.8550000000000001, 0.8999999999999999, 0.636, NaN, NaN, 0.159, 0.15600000000000003, 0.15300000000000002, 0.15600000000000003, 0.15600000000000003, 0.135, 0.168, 0.195, 0.255, 0.402, 0.42600000000000005, 0.6960000000000001, 0.777, 0.7170000000000001, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.129, 0.15600000000000003, 0.159, 0.159, 0.165, 0.14400000000000002, 0.23099999999999998, 0.399, 0.7110000000000001, 0.9570000000000001, 0.885, 0.723, 0.666, NaN, NaN, 0.15600000000000003, 0.162, 0.162, 0.168, 0.15600000000000003, 0.162, 0.17400000000000002, 0.21600000000000003, 0.27, 0.7020000000000001, 0.96, 0.45599999999999996, NaN, NaN, 0.159, 0.159, 0.162, 0.15600000000000003, 0.162, 0.135, 0.165, 0.189, 0.34800000000000003, 0.651, 0.984, 1.179, 1.197, 1.239, NaN, NaN, 0.162, 0.168, 0.162, 0.15600000000000003, 0.138, 0.162, 0.18, 0.21600000000000003, 0.342, 0.6900000000000001, 1.2480000000000002, 1.5, NaN, NaN, 0.162, 0.162, 0.15600000000000003, 0.15600000000000003, 0.162, 0.138, 0.15600000000000003, 0.168, 0.186, 0.21600000000000003, 0.24, 0.42600000000000005, 0.762, 1.182, 1.23, NaN, NaN, 0.162, 0.162, 0.15600000000000003, 0.162, 0.15600000000000003, 0.168, 0.198, 0.252, 0.396, 0.81, 1.3800000000000001, NaN, NaN, 0.159, 0.159, 0.159, 0.159, 0.159, 0.168, 0.159, 0.17700000000000002, 0.195, 0.34800000000000003, 1.1760000000000002, 1.437, 1.437, 1.446, NaN, NaN, 0.162, 0.15600000000000003, 0.162, 0.168, 0.15600000000000003, 0.162, 0.168, 0.22199999999999998, 0.43200000000000005, 0.8879999999999999, 1.3920000000000001, NaN, NaN, 0.159, 0.15300000000000002, 0.15300000000000002, 0.17700000000000002, 0.159, 0.171, 0.183, 0.23099999999999998, 0.387, 0.9930000000000001, 1.677, 1.443, 1.317, NaN, NaN, 0.159, 0.159, 0.159, 0.159, 0.159, 0.132, 0.168, 0.159, 0.28500000000000003, 0.5369999999999999, 0.6990000000000001, 1.5990000000000002, 1.293, NaN, NaN, 0.159, 0.159, 0.15300000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.171, 0.22499999999999998, 0.29100000000000004, 0.489, 0.903, 1.4489999999999998, 1.215, 1.113, NaN, NaN, 0.15600000000000003, 0.162, 0.15600000000000003, 0.162, 0.132, 0.15600000000000003, 0.17400000000000002, 0.186, 0.27, 0.5640000000000001, 0.96, 1.482, 1.158, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.165, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.138, 0.17400000000000002, 0.264, 0.5700000000000001, 1.3800000000000001, 1.5870000000000002, 1.353, 1.119, 1.056, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.162, 0.168, 0.186, 0.198, 0.252, 0.31200000000000006, 0.36, 1.0619999999999998, 1.194, NaN, NaN, 0.15600000000000003, 0.15600000000000003, 0.129, 0.15600000000000003, 0.15600000000000003, 0.15600000000000003, 0.165, 0.17400000000000002, 0.21000000000000002, 0.246, 0.30000000000000004, 0.651, 1.4969999999999999, 1.092, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.15300000000000002, 0.15300000000000002, 0.165, 0.189, 0.237, 0.261, 0.381, 0.7050000000000001, 1.365, 1.059, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.171, 0.195, 0.23099999999999998, 0.30300000000000005, 0.44099999999999995, 0.801, 1.305, 1.785, 1.0470000000000002, NaN, NaN, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.15300000000000002, 0.15300000000000002, 0.165, 0.171, 0.171, 0.22499999999999998, 0.46499999999999997, 0.9450000000000001, 1.425, 1.0410000000000001, NaN, NaN, 0.15300000000000002, 0.14700000000000002, 0.15300000000000002, 0.159, 0.15300000000000002, 0.123, 0.165, 0.165, 0.159, 0.21300000000000002, 0.201, 0.30900000000000005, 0.633, 1.305, NaN, NaN, 0.15300000000000002, 0.15600000000000003, 0.15000000000000002, 0.159, 0.15300000000000002, 0.132, 0.15600000000000003, 0.171, 0.21300000000000002, 0.243, 0.23399999999999999, 0.363, 0.663, 0.9570000000000001, 0.9059999999999999, NaN, NaN, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.126, 0.15600000000000003, 0.17700000000000002, 0.192, 0.21300000000000002, 0.276, 0.384, 0.663, 0.9690000000000001, 0.8879999999999999, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.165, 0.159, 0.15600000000000003, 0.162, 0.186, 0.23099999999999998, 0.318, 0.48, 0.777, 0.8340000000000001, 0.933, 0.8819999999999999, 0.639, NaN, NaN, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15600000000000003, 0.162, 0.183, 0.21600000000000003, 0.267, 0.321, 0.483, 0.756, 0.8280000000000001, 0.9059999999999999, 0.648, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.099, 0.15000000000000002, 0.132, 0.189, 0.21899999999999997, 0.34800000000000003, 0.34800000000000003, 0.666, 0.7080000000000001, 0.75, 0.381, NaN, NaN, 0.15000000000000002, 0.15600000000000003, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15600000000000003, 0.198, 0.24, 0.30600000000000005, 0.516, 0.516, 0.669, 0.732, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.15000000000000002, 0.129, 0.18, 0.198, 0.28200000000000003, 0.342, 0.396, 0.5489999999999999, 0.7140000000000001, 0.7080000000000001, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.159, 0.14700000000000002, 0.23099999999999998, 0.22499999999999998, 0.30000000000000004, 0.27, 0.558, 0.6120000000000001, 0.366, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.15300000000000002, 0.15600000000000003, 0.159, 0.168, 0.17400000000000002, 0.261, 0.44399999999999995, 0.777, 0.768, 0.507, 0.42300000000000004, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.165, 0.14100000000000001, 0.18, 0.189, 0.23099999999999998, 0.399, 0.5760000000000001, 0.573, 0.45599999999999996, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.159, 0.168, 0.186, 0.243, 0.45599999999999996, 0.648, 0.43799999999999994, 0.321, 0.273, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.162, 0.15000000000000002, 0.20700000000000002, 0.246, 0.252, 0.603, 0.41700000000000004, 0.384, 0.315, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.129, 0.15600000000000003, 0.159, 0.15000000000000002, 0.168, 0.23099999999999998, 0.255, 0.567, 0.672, 0.8250000000000001, 0.504, 0.34500000000000003, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14400000000000002, 0.15300000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.138, 0.189, 0.22499999999999998, 0.261, 0.399, 0.48, 0.8220000000000001, 0.654, 0.495, 0.183, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14700000000000002, 0.129, 0.15300000000000002, 0.171, 0.183, 0.246, 0.261, 0.264, 0.43499999999999994, 0.534, 0.783, 0.897, 0.44699999999999995, 0.41700000000000004, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.15600000000000003, 0.14700000000000002, 0.15300000000000002, 0.132, 0.171, 0.183, 0.21899999999999997, 0.264, 0.28500000000000003, 0.5640000000000001, 0.783, 1.0050000000000001, 0.669, 0.40800000000000003, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.11399999999999999, 0.14100000000000001, 0.14400000000000002, 0.123, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.129, 0.162, 0.183, 0.22199999999999998, 0.27, 0.42600000000000005, 0.729, 0.8310000000000001, 1.0530000000000002, 1.071, 0.5549999999999999, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15600000000000003, 0.15300000000000002, 0.129, 0.17400000000000002, 0.246, 0.366, 0.726, 0.933, 1.008, 0.9810000000000001, 0.8190000000000001, 0.801, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.171, 0.21000000000000002, 0.264, 0.43200000000000005, 0.804, 0.8610000000000001, 1.0530000000000002, 1.0619999999999998, 0.786, 0.9390000000000001, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15600000000000003, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.162, 0.189, 0.243, 0.258, 0.33, 0.6990000000000001, 0.795, 1.059, 1.0470000000000002, 0.804, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15300000000000002, 0.159, 0.171, 0.22199999999999998, 0.21300000000000002, 0.477, 0.726, 0.807, 0.9990000000000001, 0.8879999999999999, 0.8759999999999999, 0.8220000000000001, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.126, 0.126, 0.159, 0.15300000000000002, 0.171, 0.192, 0.237, 0.261, 0.321, 0.5369999999999999, 0.747, 0.639, 1.0530000000000002, 0.9450000000000001, 0.891, 0.41700000000000004, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14700000000000002, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.10200000000000001, 0.129, 0.15300000000000002, 0.159, 0.195, 0.255, 0.279, 0.333, 0.5609999999999999, 0.7050000000000001, 0.777, 1.215, 0.867, 0.885, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.123, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14700000000000002, 0.123, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.15600000000000003, 0.15600000000000003, 0.162, 0.132, 0.17700000000000002, 0.22499999999999998, 0.27, 0.276, 0.369, 0.5700000000000001, 0.6180000000000001, 0.6990000000000001, 0.8819999999999999, 1.032, 0.996, 1.077, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.15000000000000002, 0.123, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14700000000000002, 0.14400000000000002, 0.123, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.126, 0.15600000000000003, 0.159, 0.171, 0.195, 0.22799999999999998, 0.20700000000000002, 0.28800000000000003, 0.378, 0.5820000000000001, 0.72, 0.801, 0.9810000000000001, 0.972, 0.885, 1.0530000000000002, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.123, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.123, 0.123, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.12, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.15000000000000002, 0.162, 0.15300000000000002, 0.159, 0.15300000000000002, 0.159, 0.189, 0.24, 0.279, 0.33, 0.471, 0.5820000000000001, 0.645, 0.648, 0.8310000000000001, 1.0859999999999999, 1.125, 1.107, 1.173, NaN, NaN, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.11699999999999999, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.123, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.123, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14700000000000002, 0.12, 0.14700000000000002, 0.162, 0.159, 0.186, 0.237, 0.261, 0.267, 0.28500000000000003, 0.34500000000000003, 0.498, 0.627, 0.597, 0.9119999999999999, 1.014, 0.8640000000000001, 0.54, 0.336, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.15300000000000002, 0.14700000000000002, 0.14700000000000002, 0.12, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.123, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.12, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.15000000000000002, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.123, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.15300000000000002, 0.162, 0.171, 0.15600000000000003, 0.186, 0.28200000000000003, 0.29400000000000004, 0.31200000000000006, 0.336, 0.477, 0.651, 0.747, 0.8400000000000001, 0.9750000000000001, 1.158, 0.954, 0.597, 0.372, 0.28800000000000003, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14400000000000002, 0.14700000000000002, 0.099, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.099, 0.123, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.123, 0.126, 0.159, 0.165, 0.17700000000000002, 0.20700000000000002, 0.28500000000000003, 0.30000000000000004, 0.264, 0.366, 0.534, 0.7080000000000001, 0.984, 1.2120000000000002, 1.0739999999999998, 0.81, 0.54, 0.363, 0.29700000000000004, 0.201, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.123, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.168, 0.17700000000000002, 0.198, 0.237, 0.249, 0.30900000000000005, 0.336, 0.369, 0.41700000000000004, 0.5700000000000001, 0.9359999999999999, 0.9810000000000001, 1.095, 0.978, 0.6240000000000001, 0.513, 0.5369999999999999, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.12, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.129, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.15000000000000002, 0.15000000000000002, 0.162, 0.17400000000000002, 0.183, 0.21300000000000002, 0.246, 0.249, 0.318, 0.35400000000000004, 0.402, 0.46799999999999997, 0.471, 0.633, 0.8190000000000001, 1.134, 1.221, 1.0110000000000001, 0.8879999999999999, 0.7080000000000001, 0.504, 0.6060000000000001, NaN, NaN, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.12, 0.12, 0.138, 0.11399999999999999, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.093, 0.11399999999999999, 0.14400000000000002, 0.14700000000000002, 0.123, 0.15300000000000002, 0.162, 0.165, 0.18, 0.201, 0.237, 0.29700000000000004, 0.276, 0.36, 0.381, 0.46199999999999997, 0.51, 0.636, 0.8370000000000001, 0.9810000000000001, 0.672, 0.552, 0.42000000000000004, 0.48, 0.54, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14100000000000001, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.11699999999999999, 0.14100000000000001, 0.138, 0.135, 0.135, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.159, 0.132, 0.14100000000000001, 0.189, 0.21300000000000002, 0.20700000000000002, 0.22499999999999998, 0.273, 0.264, 0.42600000000000005, 0.474, 0.5700000000000001, 0.5640000000000001, 0.744, 0.984, 1.056, 0.5760000000000001, 0.43200000000000005, 0.42600000000000005, 0.336, 0.35400000000000004, 0.34800000000000003, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.12, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14700000000000002, 0.14100000000000001, 0.10800000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.12, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11699999999999999, 0.11099999999999999, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14700000000000002, 0.159, 0.171, 0.195, 0.20700000000000002, 0.23099999999999998, 0.21300000000000002, 0.255, 0.264, 0.267, 0.27, 0.28800000000000003, 0.42600000000000005, 0.7110000000000001, 0.8190000000000001, 0.642, 0.5640000000000001, 0.387, 0.369, 0.324, 0.363, 0.372, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.123, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.14400000000000002, 0.15300000000000002, 0.15600000000000003, 0.171, 0.183, 0.192, 0.186, 0.198, 0.20700000000000002, 0.23099999999999998, 0.249, 0.273, 0.261, 0.315, 0.46499999999999997, 0.5489999999999999, 0.9390000000000001, 0.891, 0.8430000000000001, 0.615, 0.369, 0.399, 0.381, 0.34500000000000003, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14700000000000002, 0.123, 0.14100000000000001, 0.11699999999999999, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.11399999999999999, 0.138, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.129, 0.168, 0.183, 0.195, 0.201, 0.20700000000000002, 0.243, 0.246, 0.23099999999999998, 0.261, 0.324, 0.369, 0.687, 0.729, 0.9239999999999999, 0.9750000000000001, 0.741, 0.387, 0.324, 0.279, 0.135, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.123, 0.123, 0.123, 0.15000000000000002, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.14400000000000002, 0.12, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14400000000000002, 0.126, 0.162, 0.17400000000000002, 0.183, 0.183, 0.195, 0.18, 0.243, 0.252, 0.24, 0.252, 0.29100000000000004, 0.387, 0.54, 0.5549999999999999, 0.681, 0.915, 0.6060000000000001, 0.5700000000000001, 0.40800000000000003, 0.29100000000000004, 0.267, 0.24, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.123, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.123, 0.11099999999999999, 0.11399999999999999, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.11399999999999999, 0.138, 0.138, 0.138, 0.12, 0.15300000000000002, 0.171, 0.189, 0.126, 0.195, 0.21300000000000002, 0.24, 0.237, 0.24, 0.273, 0.30900000000000005, 0.324, 0.44999999999999996, 0.609, 0.8580000000000001, 0.879, 0.5880000000000001, 0.366, 0.369, 0.336, 0.318, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.12, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.12, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.12, 0.11699999999999999, 0.12, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.093, 0.14400000000000002, 0.12, 0.15300000000000002, 0.171, 0.186, 0.159, 0.186, 0.195, 0.171, 0.186, 0.22799999999999998, 0.20700000000000002, 0.261, 0.28500000000000003, 0.321, 0.387, 0.8550000000000001, 0.789, 0.8370000000000001, 0.891, 0.681, 0.41700000000000004, 0.46499999999999997, 0.41100000000000003, 0.46499999999999997, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.138, 0.14700000000000002, 0.14100000000000001, 0.15000000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.12, 0.14100000000000001, 0.138, 0.14700000000000002, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.18, 0.189, 0.198, 0.192, 0.195, 0.20700000000000002, 0.22199999999999998, 0.22799999999999998, 0.246, 0.258, 0.264, 0.35700000000000004, 0.31200000000000006, 0.645, 0.9119999999999999, 0.684, 0.522, 0.41400000000000003, 0.36, 0.42000000000000004, 0.342, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14700000000000002, 0.123, 0.14700000000000002, 0.14400000000000002, 0.123, 0.14400000000000002, 0.123, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.138, 0.14400000000000002, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.14700000000000002, 0.15300000000000002, 0.159, 0.18, 0.186, 0.20400000000000001, 0.198, 0.21000000000000002, 0.22199999999999998, 0.192, 0.246, 0.273, 0.31200000000000006, 0.384, 0.42300000000000004, 0.42900000000000005, 0.759, 0.558, 0.41700000000000004, 0.29400000000000004, 0.372, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.123, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.096, 0.123, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14700000000000002, 0.15600000000000003, 0.159, 0.171, 0.18, 0.192, 0.21000000000000002, 0.201, 0.20700000000000002, 0.22499999999999998, 0.23099999999999998, 0.255, 0.28500000000000003, 0.333, 0.39, 0.45599999999999996, 0.552, 0.744, 0.46799999999999997, 0.369, 0.366, 0.34800000000000003, NaN, NaN, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.138, 0.12, 0.14100000000000001, 0.12, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11399999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.11399999999999999, 0.168, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.12, 0.17400000000000002, 0.552, 0.54, 0.546, 0.42600000000000005, 0.51, 0.48, 0.51, 0.22799999999999998, 0.20400000000000001, 0.198, 0.22199999999999998, 0.22799999999999998, 0.258, 0.27, 0.321, 0.384, 0.41700000000000004, 0.495, 0.669, 0.7080000000000001, 0.501, 0.29400000000000004, 0.27, 0.35400000000000004, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.123, 0.14400000000000002, 0.14400000000000002, 0.123, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.099, 0.12, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.11399999999999999, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.138, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.12, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.15600000000000003, 0.17400000000000002, 0.15600000000000003, 0.168, 0.201, 0.201, 0.165, 0.21600000000000003, 0.20700000000000002, 0.189, 0.23399999999999999, 0.30000000000000004, 0.318, 0.378, 0.44699999999999995, 0.41400000000000003, 0.567, 0.774, 0.7050000000000001, 0.66, 0.45299999999999996, 0.384, 0.402, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.15000000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.08700000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.165, 0.17700000000000002, 0.195, 0.192, 0.165, 0.201, 0.20700000000000002, 0.201, 0.21300000000000002, 0.21600000000000003, 0.249, 0.321, 0.42900000000000005, 0.387, 0.393, 0.399, 0.5429999999999999, 0.8490000000000001, 0.387, 0.267, 0.17700000000000002, 0.201, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.123, 0.14100000000000001, 0.14400000000000002, 0.135, 0.11699999999999999, 0.14400000000000002, 0.12, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.129, 0.17400000000000002, 0.189, 0.189, 0.17700000000000002, 0.183, 0.201, 0.20400000000000001, 0.21000000000000002, 0.21899999999999997, 0.261, 0.327, 0.43499999999999994, 0.45299999999999996, 0.5609999999999999, 0.753, 0.807, 0.41100000000000003, 0.237, 0.165, 0.14100000000000001, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.12, 0.12, 0.11699999999999999, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.11099999999999999, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.11399999999999999, 0.135, 0.138, 0.138, 0.14100000000000001, 0.15300000000000002, 0.168, 0.195, 0.22799999999999998, 0.21000000000000002, 0.21300000000000002, 0.237, 0.237, 0.21300000000000002, 0.255, 0.171, 0.5309999999999999, 0.42300000000000004, 0.5429999999999999, 0.9810000000000001, 1.0530000000000002, 0.8610000000000001, 0.8130000000000001, 0.597, 0.30300000000000005, 0.29100000000000004, 0.237, 0.22499999999999998, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.12, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.11399999999999999, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.11699999999999999, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.14400000000000002, 0.126, 0.171, 0.165, 0.198, 0.183, 0.237, 0.255, 0.276, 0.28200000000000003, 0.30000000000000004, 0.31200000000000006, 0.31200000000000006, 0.636, 0.9059999999999999, 1.0739999999999998, 1.0290000000000001, 0.765, 0.44699999999999995, 0.366, 0.29400000000000004, 0.39, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14700000000000002, 0.135, 0.14700000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.10200000000000001, 0.138, 0.11699999999999999, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.12, 0.14700000000000002, 0.162, 0.17700000000000002, 0.20400000000000001, 0.21300000000000002, 0.21899999999999997, 0.23099999999999998, 0.252, 0.243, 0.29700000000000004, 0.30900000000000005, 0.363, 0.46499999999999997, 0.9930000000000001, 0.795, 0.7110000000000001, 0.5309999999999999, 0.35100000000000003, 0.333, 0.339, 0.29700000000000004, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.132, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.138, 0.138, 0.10500000000000001, 0.138, 0.14100000000000001, 0.11399999999999999, 0.135, 0.14100000000000001, 0.138, 0.135, 0.135, 0.138, 0.14100000000000001, 0.14700000000000002, 0.15000000000000002, 0.168, 0.165, 0.198, 0.21300000000000002, 0.22499999999999998, 0.22499999999999998, 0.30000000000000004, 0.327, 0.339, 0.333, 0.381, 0.534, 0.6240000000000001, 0.9510000000000001, 0.654, 0.402, 0.342, 0.324, 0.28500000000000003, 0.267, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.12, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.14100000000000001, 0.138, 0.135, 0.138, 0.11099999999999999, 0.11699999999999999, 0.14700000000000002, 0.165, 0.186, 0.21300000000000002, 0.21300000000000002, 0.264, 0.249, 0.273, 0.28200000000000003, 0.31200000000000006, 0.378, 0.42600000000000005, 0.489, 0.633, 0.8130000000000001, 0.525, 0.41700000000000004, 0.342, 0.318, 0.267, 0.324, 0.342, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.12, 0.12, 0.14400000000000002, 0.11699999999999999, 0.138, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.09, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.162, 0.171, 0.198, 0.21899999999999997, 0.252, 0.327, 0.45299999999999996, 0.46199999999999997, 0.44099999999999995, 0.573, 0.7050000000000001, 0.732, 0.765, 0.6930000000000001, 0.43499999999999994, 0.28800000000000003, 0.33, 0.34800000000000003, 0.321, 0.387, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.138, 0.11399999999999999, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11699999999999999, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.135, 0.138, 0.14100000000000001, 0.10500000000000001, 0.135, 0.11099999999999999, 0.138, 0.135, 0.135, 0.135, 0.138, 0.14100000000000001, 0.14400000000000002, 0.15600000000000003, 0.17400000000000002, 0.195, 0.21300000000000002, 0.237, 0.276, 0.33, 0.474, 0.522, 0.5369999999999999, 0.63, 0.873, 1.095, 0.8160000000000001, 0.7140000000000001, 0.405, 0.381, 0.42000000000000004, 0.34800000000000003, 0.35400000000000004, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.12, 0.14100000000000001, 0.14400000000000002, 0.132, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.11399999999999999, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.138, 0.138, 0.135, 0.14100000000000001, 0.138, 0.069, 0.135, 0.138, 0.135, 0.138, 0.135, 0.135, 0.14100000000000001, 0.14400000000000002, 0.123, 0.15000000000000002, 0.17400000000000002, 0.186, 0.20400000000000001, 0.21899999999999997, 0.249, 0.30300000000000005, 0.29700000000000004, 0.42000000000000004, 0.498, 0.495, 0.672, 0.768, 0.972, 0.78, 0.525, 0.321, 0.324, 0.276, 0.237, 0.17400000000000002, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.135, 0.15000000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.20700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.10800000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.084, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.138, 0.135, 0.132, 0.138, 0.138, 0.14100000000000001, 0.12, 0.15300000000000002, 0.17700000000000002, 0.183, 0.20400000000000001, 0.21300000000000002, 0.24, 0.279, 0.33, 0.39, 0.363, 0.573, 0.681, 0.885, 1.0110000000000001, 0.9690000000000001, 0.369, 0.315, 0.255, 0.22499999999999998, 0.201, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.138, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.096, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.10200000000000001, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.138, 0.14100000000000001, 0.14700000000000002, 0.15600000000000003, 0.171, 0.18, 0.192, 0.20700000000000002, 0.183, 0.23399999999999999, 0.276, 0.336, 0.41400000000000003, 0.474, 0.504, 0.75, 0.966, 1.326, 1.0619999999999998, 0.5880000000000001, 0.40800000000000003, 0.342, 0.29400000000000004, 0.252, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.132, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.159, 0.171, 0.189, 0.20700000000000002, 0.23399999999999999, 0.22799999999999998, 0.237, 0.315, 0.41100000000000003, 0.501, 0.621, 0.879, 1.125, 0.9690000000000001, 0.46499999999999997, 0.42900000000000005, 0.42300000000000004, 0.393, 0.471, 0.41100000000000003, 0.405, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.135, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.138, 0.135, 0.135, 0.135, 0.11699999999999999, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.12, 0.159, 0.171, 0.183, 0.192, 0.22199999999999998, 0.243, 0.267, 0.28800000000000003, 0.339, 0.43200000000000005, 0.621, 0.8640000000000001, 1.008, 1.1760000000000002, 0.5700000000000001, 0.44999999999999996, 0.46199999999999997, 0.45599999999999996, 0.43200000000000005, 0.39, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.135, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.135, 0.138, 0.135, 0.135, 0.11099999999999999, 0.138, 0.14100000000000001, 0.14400000000000002, 0.15000000000000002, 0.165, 0.17700000000000002, 0.198, 0.21300000000000002, 0.237, 0.264, 0.29700000000000004, 0.30900000000000005, 0.35100000000000003, 0.44699999999999995, 0.5549999999999999, 0.753, 0.9750000000000001, 0.8580000000000001, 0.54, 0.5429999999999999, 0.492, 0.44399999999999995, 0.507, 0.501, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14400000000000002, 0.11699999999999999, 0.12, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.10800000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11699999999999999, 0.138, 0.138, 0.11399999999999999, 0.135, 0.11099999999999999, 0.135, 0.10800000000000001, 0.135, 0.135, 0.138, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.159, 0.162, 0.18, 0.195, 0.21300000000000002, 0.22199999999999998, 0.23399999999999999, 0.261, 0.30000000000000004, 0.342, 0.39, 0.42900000000000005, 0.495, 0.633, 0.807, 0.873, 0.648, 0.5609999999999999, 0.579, 0.5369999999999999, 0.5820000000000001, 0.54, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.11099999999999999, 0.11699999999999999, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.135, 0.093, 0.135, 0.135, 0.135, 0.10800000000000001, 0.09, 0.138, 0.14100000000000001, 0.14700000000000002, 0.135, 0.168, 0.15300000000000002, 0.171, 0.21899999999999997, 0.21000000000000002, 0.261, 0.28500000000000003, 0.315, 0.41100000000000003, 0.40800000000000003, 0.5489999999999999, 0.621, 0.759, 0.672, 0.513, 0.5880000000000001, 0.492, 0.5880000000000001, 0.63, 0.609, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.11399999999999999, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.138, 0.138, 0.135, 0.138, 0.11399999999999999, 0.135, 0.135, 0.138, 0.138, 0.14400000000000002, 0.15300000000000002, 0.14700000000000002, 0.15300000000000002, 0.165, 0.18, 0.23399999999999999, 0.22499999999999998, 0.23099999999999998, 0.21300000000000002, 0.28800000000000003, 0.36, 0.40800000000000003, 0.45899999999999996, 0.45899999999999996, 0.5760000000000001, 0.633, 0.771, 0.642, 0.663, 0.597, 0.687, 0.567, 0.363, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.135, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.138, 0.11699999999999999, 0.11099999999999999, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.14100000000000001, 0.14400000000000002, 0.15300000000000002, 0.168, 0.189, 0.21000000000000002, 0.243, 0.258, 0.315, 0.35700000000000004, 0.381, 0.43799999999999994, 0.504, 0.642, 0.756, 0.7110000000000001, 0.678, 0.6240000000000001, 0.45299999999999996, 0.35700000000000004, 0.28500000000000003, 0.28200000000000003, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.12, 0.096, 0.14400000000000002, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.12, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.135, 0.138, 0.093, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.11399999999999999, 0.138, 0.135, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.138, 0.135, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.17700000000000002, 0.192, 0.21300000000000002, 0.23399999999999999, 0.21600000000000003, 0.27, 0.276, 0.28200000000000003, 0.273, 0.29700000000000004, 0.35100000000000003, 0.528, 0.63, 0.9239999999999999, 0.8939999999999999, 0.9299999999999999, 0.654, 0.501, 0.27, 0.27, 0.30300000000000005, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.11399999999999999, 0.11699999999999999, 0.11099999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.11699999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.11399999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.10200000000000001, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.138, 0.138, 0.132, 0.14400000000000002, 0.11099999999999999, 0.138, 0.14100000000000001, 0.14700000000000002, 0.165, 0.17700000000000002, 0.198, 0.186, 0.261, 0.279, 0.29700000000000004, 0.327, 0.258, 0.333, 0.486, 0.678, 0.7140000000000001, 0.903, 0.9450000000000001, 0.804, 0.7140000000000001, 0.6240000000000001, 0.522, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.132, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.10500000000000001, 0.11399999999999999, 0.135, 0.135, 0.135, 0.10200000000000001, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.10500000000000001, 0.138, 0.14100000000000001, 0.138, 0.14400000000000002, 0.15300000000000002, 0.17400000000000002, 0.21899999999999997, 0.21000000000000002, 0.35400000000000004, 0.273, 0.42000000000000004, 0.486, 0.678, 0.915, 0.9870000000000001, 0.9359999999999999, 0.915, 0.8819999999999999, 0.9390000000000001, 0.903, 0.927, 0.9690000000000001, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.132, 0.132, 0.11399999999999999, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.10500000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.135, 0.138, 0.10800000000000001, 0.138, 0.138, 0.11099999999999999, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.138, 0.11099999999999999, 0.14700000000000002, 0.162, 0.21600000000000003, 0.237, 0.246, 0.264, 0.29100000000000004, 0.405, 0.498, 0.5700000000000001, 0.615, 0.738, 0.873, 0.795, 0.948, 0.909, 0.753, 0.921, 0.774, 0.879, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.132, 0.11399999999999999, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14700000000000002, 0.11399999999999999, 0.138, 0.135, 0.138, 0.11699999999999999, 0.11699999999999999, 0.10200000000000001, 0.10800000000000001, 0.11399999999999999, 0.138, 0.135, 0.135, 0.132, 0.132, 0.11399999999999999, 0.135, 0.132, 0.135, 0.11399999999999999, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.15000000000000002, 0.159, 0.21899999999999997, 0.267, 0.318, 0.342, 0.44099999999999995, 0.5549999999999999, 0.72, 0.99, 0.948, 0.996, 0.948, 0.9359999999999999, 0.9690000000000001, 0.9990000000000001, 0.801, 0.498, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.135, 0.14100000000000001, 0.135, 0.14100000000000001, 0.14100000000000001, 0.138, 0.135, 0.135, 0.135, 0.10800000000000001, 0.138, 0.10800000000000001, 0.135, 0.11399999999999999, 0.132, 0.135, 0.135, 0.135, 0.138, 0.14100000000000001, 0.14400000000000002, 0.129, 0.15600000000000003, 0.165, 0.18, 0.189, 0.29700000000000004, 0.324, 0.36, 0.51, 0.663, 0.879, 0.9239999999999999, 0.8999999999999999, 0.78, 0.8999999999999999, 0.909, 0.732, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.11399999999999999, 0.135, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.10800000000000001, 0.138, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.138, 0.132, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11399999999999999, 0.138, 0.14400000000000002, 0.14400000000000002, 0.132, 0.165, 0.171, 0.186, 0.20700000000000002, 0.23099999999999998, 0.249, 0.279, 0.339, 0.396, 0.41400000000000003, 0.528, 0.984, 0.978, 0.972, 0.8340000000000001, 0.9179999999999999, 0.9299999999999999, 1.1400000000000001, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.135, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.11099999999999999, 0.138, 0.11099999999999999, 0.10200000000000001, 0.10800000000000001, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11399999999999999, 0.132, 0.135, 0.138, 0.138, 0.135, 0.14100000000000001, 0.14400000000000002, 0.15600000000000003, 0.162, 0.138, 0.168, 0.18, 0.201, 0.22499999999999998, 0.261, 0.28500000000000003, 0.30600000000000005, 0.35700000000000004, 0.45299999999999996, 0.759, 0.9570000000000001, 1.05, 0.954, 0.747, 0.738, 0.573, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.138, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.11399999999999999, 0.138, 0.135, 0.138, 0.138, 0.135, 0.135, 0.138, 0.10200000000000001, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.11399999999999999, 0.138, 0.138, 0.138, 0.14100000000000001, 0.15000000000000002, 0.165, 0.15300000000000002, 0.18, 0.201, 0.22499999999999998, 0.237, 0.264, 0.30000000000000004, 0.363, 0.405, 0.579, 1.0470000000000002, 0.9870000000000001, 0.867, 0.489, 0.363, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.138, 0.11699999999999999, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.10500000000000001, 0.135, 0.135, 0.11099999999999999, 0.138, 0.138, 0.132, 0.093, 0.10200000000000001, 0.135, 0.135, 0.135, 0.10500000000000001, 0.135, 0.132, 0.135, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.11399999999999999, 0.138, 0.138, 0.11699999999999999, 0.14700000000000002, 0.14700000000000002, 0.171, 0.192, 0.20400000000000001, 0.21300000000000002, 0.21600000000000003, 0.243, 0.264, 0.29700000000000004, 0.35100000000000003, 0.42900000000000005, 0.5549999999999999, 1.215, 1.185, 1.311, 1.107, 0.8430000000000001, 0.513, 0.41700000000000004, 0.333, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.069, 0.138, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.11099999999999999, 0.11699999999999999, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.165, 0.17700000000000002, 0.198, 0.22199999999999998, 0.249, 0.252, 0.267, 0.30300000000000005, 0.30300000000000005, 0.513, 0.675, 1.251, 1.125, 1.131, 0.9870000000000001, 0.7110000000000001, 0.639, 0.603, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.14100000000000001, 0.11099999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.135, 0.138, 0.138, 0.138, 0.138, 0.135, 0.135, 0.138, 0.135, 0.10500000000000001, 0.135, 0.138, 0.11399999999999999, 0.10800000000000001, 0.11399999999999999, 0.10800000000000001, 0.135, 0.11099999999999999, 0.132, 0.135, 0.135, 0.11399999999999999, 0.14100000000000001, 0.14400000000000002, 0.15300000000000002, 0.168, 0.159, 0.198, 0.22499999999999998, 0.255, 0.23399999999999999, 0.31200000000000006, 0.40800000000000003, 0.54, 0.6060000000000001, 0.5940000000000001, 0.996, 1.08, 0.96, 0.9059999999999999, 0.8160000000000001, 0.768, 0.678, 0.744, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.12, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.138, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11099999999999999, 0.138, 0.10200000000000001, 0.132, 0.132, 0.135, 0.138, 0.11699999999999999, 0.123, 0.15300000000000002, 0.162, 0.186, 0.20400000000000001, 0.22199999999999998, 0.237, 0.279, 0.35400000000000004, 0.44999999999999996, 0.6960000000000001, 0.891, 0.921, 0.735, 0.723, 0.687, 0.666, 0.522, 0.6060000000000001, 0.663, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.12, 0.12, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.132, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.138, 0.138, 0.11699999999999999, 0.135, 0.138, 0.138, 0.132, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.11399999999999999, 0.14100000000000001, 0.15000000000000002, 0.168, 0.14400000000000002, 0.195, 0.21300000000000002, 0.243, 0.249, 0.30900000000000005, 0.366, 0.43200000000000005, 0.63, 0.948, 0.801, 0.609, 0.591, 0.5609999999999999, 0.5700000000000001, 0.558, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.135, 0.138, 0.135, 0.132, 0.11399999999999999, 0.138, 0.11399999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.138, 0.14400000000000002, 0.14700000000000002, 0.162, 0.17400000000000002, 0.192, 0.20700000000000002, 0.255, 0.28200000000000003, 0.28800000000000003, 0.35700000000000004, 0.44099999999999995, 0.627, 1.0110000000000001, 0.621, 0.609, 0.573, 0.519, 0.513, 0.41100000000000003, 0.363, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.11099999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.07200000000000001, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.138, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.11399999999999999, 0.135, 0.132, 0.132, 0.135, 0.135, 0.10500000000000001, 0.10800000000000001, 0.135, 0.138, 0.14700000000000002, 0.159, 0.162, 0.18, 0.20700000000000002, 0.21899999999999997, 0.246, 0.30900000000000005, 0.34800000000000003, 0.44099999999999995, 0.5609999999999999, 0.8879999999999999, 0.765, 0.639, 0.42000000000000004, 0.45599999999999996, 0.489, 0.372, 0.387, 0.34800000000000003, NaN, NaN, 0.14100000000000001, 0.135, 0.11099999999999999, 0.138, 0.11099999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.10800000000000001, 0.138, 0.09, 0.135, 0.14100000000000001, 0.138, 0.11099999999999999, 0.138, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.138, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.138, 0.14400000000000002, 0.15000000000000002, 0.159, 0.17400000000000002, 0.198, 0.23399999999999999, 0.261, 0.279, 0.276, 0.276, 0.48, 0.636, 0.8250000000000001, 1.482, 0.573, 0.43799999999999994, 0.393, 0.35700000000000004, 0.34800000000000003, 0.267, 0.22199999999999998, 0.22199999999999998, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.138, 0.123, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.135, 0.138, 0.10500000000000001, 0.138, 0.138, 0.138, 0.135, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.11399999999999999, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.135, 0.135, 0.132, 0.14100000000000001, 0.14100000000000001, 0.15000000000000002, 0.171, 0.18, 0.195, 0.22199999999999998, 0.252, 0.34500000000000003, 0.405, 0.573, 0.741, 0.8490000000000001, 0.507, 0.369, 0.29400000000000004, 0.243, 0.20400000000000001, 0.17700000000000002, 0.138, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.135, 0.135, 0.14400000000000002, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.11399999999999999, 0.138, 0.138, 0.14100000000000001, 0.138, 0.135, 0.138, 0.138, 0.135, 0.135, 0.138, 0.135, 0.10800000000000001, 0.135, 0.10800000000000001, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.138, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.162, 0.183, 0.20700000000000002, 0.24, 0.29400000000000004, 0.333, 0.45899999999999996, 0.525, 0.8430000000000001, 0.8130000000000001, 0.369, 0.28500000000000003, 0.23099999999999998, 0.189, 0.171, 0.159, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.10500000000000001, 0.14400000000000002, 0.14400000000000002, 0.10800000000000001, 0.135, 0.11399999999999999, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.138, 0.11099999999999999, 0.138, 0.138, 0.135, 0.135, 0.135, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.135, 0.138, 0.14100000000000001, 0.126, 0.159, 0.165, 0.189, 0.22499999999999998, 0.246, 0.339, 0.387, 0.513, 0.765, 0.948, 0.678, 0.321, 0.30000000000000004, 0.252, 0.195, 0.21600000000000003, 0.186, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.12, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.12, 0.11399999999999999, 0.14100000000000001, 0.135, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11099999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.138, 0.10800000000000001, 0.138, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.129, 0.132, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.14100000000000001, 0.15000000000000002, 0.159, 0.17400000000000002, 0.171, 0.21600000000000003, 0.28500000000000003, 0.372, 0.507, 0.732, 1.056, 0.5640000000000001, 0.36, 0.315, 0.30300000000000005, 0.273, 0.23399999999999999, 0.321, 0.28500000000000003, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.11699999999999999, 0.11399999999999999, 0.138, 0.132, 0.129, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.138, 0.135, 0.138, 0.135, 0.138, 0.132, 0.135, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.138, 0.138, 0.14400000000000002, 0.15600000000000003, 0.168, 0.195, 0.22199999999999998, 0.30300000000000005, 0.36, 0.579, 0.8550000000000001, 1.077, 0.501, 0.339, 0.327, 0.30300000000000005, 0.255, 0.27, NaN, NaN, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.132, 0.11099999999999999, 0.14400000000000002, 0.138, 0.138, 0.14100000000000001, 0.138, 0.11399999999999999, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.132, 0.135, 0.11399999999999999, 0.135, 0.10800000000000001, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.135, 0.11699999999999999, 0.14700000000000002, 0.15300000000000002, 0.183, 0.21000000000000002, 0.21000000000000002, 0.246, 0.315, 0.39, 0.558, 0.768, 0.909, 0.6180000000000001, 0.29400000000000004, 0.27, 0.276, 0.276, 0.276, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.135, 0.138, 0.132, 0.138, 0.11399999999999999, 0.11699999999999999, 0.138, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.11399999999999999, 0.11399999999999999, 0.11699999999999999, 0.138, 0.138, 0.135, 0.132, 0.132, 0.132, 0.135, 0.099, 0.11099999999999999, 0.132, 0.132, 0.10500000000000001, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.10800000000000001, 0.14100000000000001, 0.126, 0.162, 0.192, 0.237, 0.273, 0.321, 0.399, 0.513, 0.657, 0.795, 1.083, 0.585, 0.29100000000000004, 0.273, 0.28500000000000003, 0.267, 0.22499999999999998, 0.321, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.135, 0.129, 0.11099999999999999, 0.138, 0.138, 0.138, 0.11399999999999999, 0.138, 0.135, 0.14100000000000001, 0.135, 0.138, 0.135, 0.135, 0.138, 0.10800000000000001, 0.138, 0.132, 0.135, 0.132, 0.135, 0.138, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.10500000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.14100000000000001, 0.15300000000000002, 0.18, 0.201, 0.22799999999999998, 0.267, 0.29400000000000004, 0.369, 0.519, 0.627, 0.8490000000000001, 1.0290000000000001, 0.915, 0.29700000000000004, 0.273, 0.22499999999999998, 0.30300000000000005, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.138, 0.11699999999999999, 0.135, 0.132, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.135, 0.138, 0.138, 0.11099999999999999, 0.138, 0.135, 0.138, 0.135, 0.138, 0.132, 0.135, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.135, 0.135, 0.14100000000000001, 0.15000000000000002, 0.189, 0.261, 0.35100000000000003, 0.42000000000000004, 0.495, 0.735, 0.9810000000000001, 1.113, 0.45299999999999996, 0.261, 0.267, 0.249, 0.255, 0.273, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.126, 0.135, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.135, 0.11399999999999999, 0.135, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.138, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.11399999999999999, 0.138, 0.14700000000000002, 0.165, 0.20700000000000002, 0.237, 0.29700000000000004, 0.327, 0.375, 0.44099999999999995, 0.741, 0.927, 0.8430000000000001, 0.30900000000000005, 0.23099999999999998, 0.20700000000000002, 0.17700000000000002, 0.165, 0.10500000000000001, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.135, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.135, 0.11399999999999999, 0.138, 0.135, 0.11399999999999999, 0.135, 0.099, 0.135, 0.132, 0.10200000000000001, 0.135, 0.135, 0.11099999999999999, 0.135, 0.10500000000000001, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.135, 0.132, 0.135, 0.138, 0.14400000000000002, 0.14700000000000002, 0.15600000000000003, 0.186, 0.246, 0.30300000000000005, 0.339, 0.396, 0.5489999999999999, 0.663, 0.8819999999999999, 0.5640000000000001, 0.255, 0.21600000000000003, 0.201, 0.18, 0.162, 0.162, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.135, 0.129, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.135, 0.138, 0.138, 0.14100000000000001, 0.135, 0.138, 0.10800000000000001, 0.135, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10500000000000001, 0.14100000000000001, 0.15000000000000002, 0.17700000000000002, 0.168, 0.22199999999999998, 0.249, 0.261, 0.35100000000000003, 0.387, 0.513, 0.759, 1.0410000000000001, 0.651, 0.35100000000000003, 0.333, 0.267, 0.195, 0.21899999999999997, 0.201, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.138, 0.14100000000000001, 0.138, 0.135, 0.138, 0.138, 0.135, 0.132, 0.11399999999999999, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10500000000000001, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11399999999999999, 0.14100000000000001, 0.15000000000000002, 0.162, 0.162, 0.189, 0.21899999999999997, 0.264, 0.29700000000000004, 0.30000000000000004, 0.279, 0.375, 0.489, 0.597, 0.8130000000000001, 1.0530000000000002, 0.5489999999999999, 0.41700000000000004, 0.339, 0.327, 0.315, 0.339, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.14100000000000001, 0.135, 0.132, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.135, 0.135, 0.135, 0.135, 0.10200000000000001, 0.135, 0.135, 0.135, 0.10800000000000001, 0.132, 0.132, 0.135, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.138, 0.138, 0.11399999999999999, 0.15000000000000002, 0.15600000000000003, 0.168, 0.201, 0.21899999999999997, 0.237, 0.261, 0.31200000000000006, 0.43499999999999994, 0.591, 0.9390000000000001, 0.732, 0.609, 0.483, 0.363, 0.315, 0.30900000000000005, 0.22199999999999998, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.135, 0.138, 0.138, 0.138, 0.14100000000000001, 0.135, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.093, 0.138, 0.138, 0.135, 0.135, 0.11099999999999999, 0.135, 0.138, 0.132, 0.135, 0.132, 0.11399999999999999, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.14100000000000001, 0.14700000000000002, 0.162, 0.18, 0.186, 0.20700000000000002, 0.255, 0.279, 0.387, 0.42900000000000005, 0.573, 1.191, 0.807, 0.5609999999999999, 0.375, 0.339, 0.315, 0.30300000000000005, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.135, 0.129, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.10200000000000001, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.11399999999999999, 0.135, 0.10500000000000001, 0.135, 0.11099999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.14100000000000001, 0.138, 0.14100000000000001, 0.15000000000000002, 0.15000000000000002, 0.159, 0.18, 0.195, 0.22499999999999998, 0.267, 0.30000000000000004, 0.35100000000000003, 0.46799999999999997, 0.558, 0.6960000000000001, 0.723, 0.774, 0.672, 0.477, 0.30000000000000004, 0.30000000000000004, 0.249, 0.276, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11399999999999999, 0.14100000000000001, 0.138, 0.135, 0.138, 0.14100000000000001, 0.138, 0.132, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11399999999999999, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.135, 0.138, 0.135, 0.10800000000000001, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.138, 0.135, 0.12, 0.159, 0.17700000000000002, 0.189, 0.23399999999999999, 0.276, 0.315, 0.35100000000000003, 0.43499999999999994, 0.5609999999999999, 0.738, 0.7020000000000001, 0.726, 0.528, 0.363, 0.31200000000000006, 0.324, 0.31200000000000006, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.138, 0.10800000000000001, 0.11399999999999999, 0.14100000000000001, 0.138, 0.138, 0.138, 0.10500000000000001, 0.10800000000000001, 0.138, 0.129, 0.138, 0.12, 0.138, 0.138, 0.14100000000000001, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.129, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.135, 0.138, 0.14700000000000002, 0.15000000000000002, 0.165, 0.189, 0.192, 0.22199999999999998, 0.252, 0.29700000000000004, 0.381, 0.44399999999999995, 0.5820000000000001, 0.8220000000000001, 0.639, 0.339, 0.24, 0.258, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.135, 0.10800000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.135, 0.14100000000000001, 0.138, 0.11399999999999999, 0.138, 0.135, 0.135, 0.138, 0.135, 0.132, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.10800000000000001, 0.135, 0.132, 0.138, 0.12, 0.14700000000000002, 0.162, 0.171, 0.17700000000000002, 0.195, 0.20700000000000002, 0.318, 0.339, 0.5369999999999999, 0.684, 0.8759999999999999, 0.8400000000000001, 0.678, 0.5640000000000001, 0.324, 0.21600000000000003, 0.22799999999999998, 0.189, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.08700000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.129, 0.135, 0.14100000000000001, 0.138, 0.138, 0.10800000000000001, 0.138, 0.135, 0.138, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.135, 0.12, 0.15000000000000002, 0.162, 0.171, 0.198, 0.243, 0.27, 0.29400000000000004, 0.384, 0.5309999999999999, 0.744, 0.9119999999999999, 0.8250000000000001, 0.645, 0.492, 0.378, 0.342, 0.267, 0.23099999999999998, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11099999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.11699999999999999, 0.138, 0.135, 0.138, 0.135, 0.135, 0.138, 0.138, 0.135, 0.135, 0.138, 0.135, 0.10200000000000001, 0.132, 0.132, 0.132, 0.132, 0.11399999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.14100000000000001, 0.14400000000000002, 0.15600000000000003, 0.168, 0.15600000000000003, 0.21000000000000002, 0.279, 0.396, 0.471, 0.585, 0.909, 0.9239999999999999, 0.909, 0.867, 0.6240000000000001, 0.513, 0.41400000000000003, 0.378, 0.276, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14400000000000002, 0.11099999999999999, 0.138, 0.09, 0.14100000000000001, 0.138, 0.135, 0.138, 0.138, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.132, 0.135, 0.10800000000000001, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.135, 0.132, 0.132, 0.135, 0.138, 0.15600000000000003, 0.14400000000000002, 0.20700000000000002, 0.22799999999999998, 0.318, 0.42000000000000004, 0.639, 0.9059999999999999, 1.068, 1.1400000000000001, 0.8939999999999999, 0.46199999999999997, 0.41400000000000003, 0.396, 0.40800000000000003, 0.402, 0.396, 0.40800000000000003, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11399999999999999, 0.14100000000000001, 0.11699999999999999, 0.135, 0.138, 0.138, 0.093, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.138, 0.135, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.129, 0.11099999999999999, 0.11099999999999999, 0.138, 0.14700000000000002, 0.168, 0.17400000000000002, 0.189, 0.21300000000000002, 0.29400000000000004, 0.36, 0.471, 0.6060000000000001, 0.726, 0.9570000000000001, 1.1400000000000001, 1.113, 0.777, 0.405, 0.396, 0.381, 0.39, 0.315, 0.372, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.11399999999999999, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.11099999999999999, 0.135, 0.138, 0.14100000000000001, 0.138, 0.135, 0.138, 0.138, 0.135, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10500000000000001, 0.138, 0.15600000000000003, 0.165, 0.18, 0.20700000000000002, 0.237, 0.387, 0.558, 0.7050000000000001, 0.771, 1.05, 0.8490000000000001, 0.45899999999999996, 0.30900000000000005, 0.30300000000000005, 0.315, 0.30300000000000005, 0.29700000000000004, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11099999999999999, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.135, 0.135, 0.132, 0.138, 0.138, 0.11399999999999999, 0.138, 0.138, 0.138, 0.11399999999999999, 0.10800000000000001, 0.138, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.129, 0.135, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.135, 0.129, 0.132, 0.132, 0.132, 0.129, 0.138, 0.132, 0.135, 0.138, 0.15300000000000002, 0.162, 0.168, 0.186, 0.21300000000000002, 0.267, 0.342, 0.381, 0.44099999999999995, 0.7050000000000001, 0.8640000000000001, 0.609, 0.507, 0.504, 0.45599999999999996, 0.384, 0.29700000000000004, 0.29400000000000004, 0.29400000000000004, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.138, 0.11399999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.11099999999999999, 0.138, 0.11399999999999999, 0.138, 0.135, 0.135, 0.135, 0.129, 0.138, 0.138, 0.135, 0.138, 0.093, 0.135, 0.135, 0.132, 0.138, 0.10200000000000001, 0.135, 0.132, 0.132, 0.10500000000000001, 0.132, 0.10500000000000001, 0.132, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.135, 0.081, 0.14400000000000002, 0.15600000000000003, 0.159, 0.195, 0.21600000000000003, 0.28200000000000003, 0.28200000000000003, 0.35400000000000004, 0.45299999999999996, 0.741, 0.867, 0.792, 0.42000000000000004, 0.471, 0.46499999999999997, 0.45899999999999996, 0.45299999999999996, 0.44099999999999995, 0.43799999999999994, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.135, 0.14100000000000001, 0.138, 0.14400000000000002, 0.129, 0.135, 0.135, 0.138, 0.138, 0.138, 0.138, 0.135, 0.081, 0.11099999999999999, 0.132, 0.135, 0.135, 0.11099999999999999, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.135, 0.132, 0.135, 0.14700000000000002, 0.14400000000000002, 0.165, 0.171, 0.195, 0.22799999999999998, 0.237, 0.30900000000000005, 0.399, 0.44699999999999995, 0.663, 0.9059999999999999, 0.6900000000000001, 0.46199999999999997, 0.44699999999999995, 0.42000000000000004, 0.396, 0.36, 0.29400000000000004, 0.198, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.11699999999999999, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.11099999999999999, 0.138, 0.135, 0.138, 0.135, 0.132, 0.138, 0.135, 0.138, 0.14100000000000001, 0.138, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.138, 0.14700000000000002, 0.15000000000000002, 0.17700000000000002, 0.201, 0.21600000000000003, 0.21899999999999997, 0.22199999999999998, 0.28200000000000003, 0.339, 0.43499999999999994, 0.669, 0.885, 0.879, 0.744, 0.45899999999999996, 0.29700000000000004, 0.21899999999999997, 0.198, 0.17700000000000002, 0.165, 0.15000000000000002, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.135, 0.135, 0.138, 0.135, 0.132, 0.138, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.138, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.12, 0.14700000000000002, 0.15600000000000003, 0.17700000000000002, 0.21000000000000002, 0.198, 0.21000000000000002, 0.237, 0.24, 0.363, 0.5820000000000001, 0.9119999999999999, 0.921, 0.9810000000000001, 0.9930000000000001, 0.5309999999999999, 0.315, 0.23099999999999998, 0.189, 0.165, 0.135, NaN, NaN, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.135, 0.138, 0.129, 0.11399999999999999, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.138, 0.15300000000000002, 0.15300000000000002, 0.17700000000000002, 0.23099999999999998, 0.255, 0.264, 0.318, 0.366, 0.45899999999999996, 0.8250000000000001, 1.008, 0.915, 0.45899999999999996, 0.43799999999999994, 0.363, 0.273, 0.21600000000000003, 0.198, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.135, 0.11099999999999999, 0.138, 0.138, 0.14100000000000001, 0.129, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.135, 0.138, 0.10200000000000001, 0.10200000000000001, 0.10800000000000001, 0.14100000000000001, 0.138, 0.11099999999999999, 0.135, 0.135, 0.132, 0.135, 0.132, 0.09, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.135, 0.138, 0.14400000000000002, 0.15600000000000003, 0.18, 0.22799999999999998, 0.255, 0.321, 0.327, 0.42000000000000004, 0.522, 0.633, 0.768, 1.0170000000000001, 0.81, 0.6960000000000001, 0.609, 0.45299999999999996, 0.324, 0.29400000000000004, 0.28200000000000003, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.11099999999999999, 0.14100000000000001, 0.135, 0.135, 0.138, 0.135, 0.129, 0.10800000000000001, 0.132, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.14100000000000001, 0.14400000000000002, 0.132, 0.168, 0.159, 0.27, 0.363, 0.41100000000000003, 0.44099999999999995, 0.5820000000000001, 0.8400000000000001, 0.909, 0.756, 0.6900000000000001, 0.387, 0.477, 0.342, 0.30000000000000004, 0.29100000000000004, 0.29100000000000004, NaN, NaN, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.11699999999999999, 0.11399999999999999, 0.11099999999999999, 0.138, 0.138, 0.138, 0.135, 0.11099999999999999, 0.135, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.138, 0.132, 0.135, 0.138, 0.132, 0.132, 0.138, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.11399999999999999, 0.11099999999999999, 0.135, 0.14100000000000001, 0.15000000000000002, 0.159, 0.168, 0.195, 0.186, 0.252, 0.324, 0.498, 0.72, 0.9359999999999999, 0.942, 0.522, 0.474, 0.276, 0.318, 0.336, 0.30000000000000004, NaN, NaN, 0.138, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.135, 0.138, 0.11399999999999999, 0.138, 0.129, 0.11699999999999999, 0.11699999999999999, 0.138, 0.11699999999999999, 0.138, 0.135, 0.138, 0.10800000000000001, 0.138, 0.135, 0.135, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11399999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.138, 0.14100000000000001, 0.15000000000000002, 0.15300000000000002, 0.168, 0.123, 0.20400000000000001, 0.23399999999999999, 0.267, 0.30900000000000005, 0.387, 0.501, 0.6240000000000001, 0.954, 1.0170000000000001, 0.678, 0.633, 0.483, 0.36, 0.21300000000000002, 0.22799999999999998, NaN, NaN, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.132, 0.129, 0.11699999999999999, 0.14100000000000001, 0.138, 0.135, 0.138, 0.11099999999999999, 0.135, 0.138, 0.138, 0.135, 0.132, 0.135, 0.10800000000000001, 0.11399999999999999, 0.138, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.135, 0.129, 0.129, 0.135, 0.129, 0.135, 0.11099999999999999, 0.14100000000000001, 0.14700000000000002, 0.165, 0.171, 0.171, 0.249, 0.28500000000000003, 0.30900000000000005, 0.375, 0.501, 0.753, 1.203, 1.0350000000000001, 0.765, 0.54, 0.495, 0.384, 0.327, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.11699999999999999, 0.138, 0.138, 0.138, 0.14100000000000001, 0.14100000000000001, 0.11099999999999999, 0.14100000000000001, 0.138, 0.135, 0.11099999999999999, 0.129, 0.138, 0.138, 0.138, 0.135, 0.11099999999999999, 0.11699999999999999, 0.138, 0.138, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.10500000000000001, 0.135, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.135, 0.138, 0.14400000000000002, 0.129, 0.192, 0.21300000000000002, 0.24, 0.28500000000000003, 0.33, 0.501, 0.513, 0.753, 1.149, 0.579, 0.5549999999999999, 0.43499999999999994, 0.261, 0.171, 0.183, NaN, NaN, 0.14400000000000002, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.051000000000000004, 0.138, 0.138, 0.138, 0.135, 0.138, 0.084, 0.138, 0.138, 0.138, 0.135, 0.138, 0.129, 0.14100000000000001, 0.138, 0.138, 0.138, 0.14100000000000001, 0.135, 0.14100000000000001, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.135, 0.132, 0.132, 0.14100000000000001, 0.138, 0.14400000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.20400000000000001, 0.23399999999999999, 0.24, 0.28200000000000003, 0.34800000000000003, 0.43200000000000005, 0.5700000000000001, 0.8400000000000001, 0.972, 1.0979999999999999, 0.54, 0.30600000000000005, 0.24, 0.186, 0.138, 0.15000000000000002, NaN, NaN, 0.14100000000000001, 0.135, 0.135, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.10800000000000001, 0.138, 0.132, 0.135, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.14700000000000002, 0.132, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.135, 0.135, 0.11099999999999999, 0.15000000000000002, 0.165, 0.192, 0.22199999999999998, 0.276, 0.30600000000000005, 0.384, 0.51, 0.663, 1.137, 0.573, 0.375, 0.261, 0.20700000000000002, 0.17700000000000002, 0.159, NaN, NaN, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.11099999999999999, 0.138, 0.138, 0.135, 0.135, 0.11399999999999999, 0.132, 0.132, 0.135, 0.11699999999999999, 0.135, 0.138, 0.135, 0.135, 0.138, 0.10200000000000001, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.135, 0.129, 0.132, 0.129, 0.135, 0.135, 0.135, 0.14400000000000002, 0.15300000000000002, 0.17400000000000002, 0.192, 0.237, 0.276, 0.324, 0.42900000000000005, 0.507, 0.723, 1.182, 1.02, 1.254, 0.363, 0.318, 0.30000000000000004, 0.28200000000000003, 0.237, 0.246, 0.237, NaN, NaN, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.132, 0.129, 0.138, 0.135, 0.138, 0.135, 0.135, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.10500000000000001, 0.135, 0.11099999999999999, 0.135, 0.135, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.15000000000000002, 0.135, 0.14400000000000002, 0.15000000000000002, 0.17700000000000002, 0.195, 0.261, 0.30600000000000005, 0.339, 0.43499999999999994, 0.585, 0.735, 1.0470000000000002, 0.603, 0.30300000000000005, 0.273, 0.279, 0.261, 0.258, 0.24, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.138, 0.135, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.11399999999999999, 0.138, 0.135, 0.135, 0.129, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11399999999999999, 0.14100000000000001, 0.135, 0.10800000000000001, 0.132, 0.135, 0.11099999999999999, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.11099999999999999, 0.10800000000000001, 0.132, 0.138, 0.14400000000000002, 0.15600000000000003, 0.165, 0.20700000000000002, 0.24, 0.237, 0.321, 0.35100000000000003, 0.43799999999999994, 0.684, 0.8699999999999999, 0.372, 0.23399999999999999, 0.29400000000000004, 0.246, 0.252, 0.23399999999999999, 0.22799999999999998, NaN, NaN, 0.138, 0.138, 0.138, 0.135, 0.14100000000000001, 0.14100000000000001, 0.135, 0.135, 0.132, 0.129, 0.138, 0.138, 0.135, 0.138, 0.132, 0.138, 0.132, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.135, 0.129, 0.129, 0.135, 0.129, 0.135, 0.129, 0.11099999999999999, 0.14100000000000001, 0.15300000000000002, 0.135, 0.20700000000000002, 0.279, 0.35700000000000004, 0.41100000000000003, 0.471, 0.603, 0.927, 0.42900000000000005, 0.264, 0.22799999999999998, 0.21600000000000003, 0.183, 0.21600000000000003, NaN, NaN, 0.138, 0.138, 0.135, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.135, 0.135, 0.135, 0.126, 0.135, 0.11699999999999999, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10500000000000001, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10500000000000001, 0.129, 0.09, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.15300000000000002, 0.132, 0.132, 0.11099999999999999, 0.14100000000000001, 0.15600000000000003, 0.14400000000000002, 0.20700000000000002, 0.237, 0.321, 0.41700000000000004, 0.615, 0.96, 0.753, 0.381, 0.28800000000000003, 0.255, 0.23099999999999998, 0.23099999999999998, 0.24, 0.237, NaN, NaN, 0.138, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.138, 0.129, 0.138, 0.135, 0.14100000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.10500000000000001, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10500000000000001, 0.132, 0.14100000000000001, 0.14400000000000002, 0.20400000000000001, 0.264, 0.33, 0.43200000000000005, 0.474, 0.744, 0.954, 0.96, 0.5760000000000001, 0.372, 0.30600000000000005, 0.258, 0.24, 0.198, 0.24, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.138, 0.138, 0.135, 0.132, 0.138, 0.126, 0.126, 0.10800000000000001, 0.138, 0.135, 0.132, 0.135, 0.135, 0.132, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.14100000000000001, 0.10800000000000001, 0.129, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.10800000000000001, 0.11099999999999999, 0.14100000000000001, 0.168, 0.21000000000000002, 0.264, 0.333, 0.396, 0.5549999999999999, 0.726, 0.978, 0.684, 0.405, 0.22499999999999998, 0.237, 0.22199999999999998, 0.20400000000000001, 0.18, NaN, NaN, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.09, 0.135, 0.132, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.14100000000000001, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.14100000000000001, 0.132, 0.135, 0.135, 0.132, 0.135, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.15000000000000002, 0.17700000000000002, 0.21300000000000002, 0.261, 0.35400000000000004, 0.498, 0.672, 0.792, 0.8160000000000001, 0.30600000000000005, 0.20400000000000001, 0.17400000000000002, 0.162, 0.15600000000000003, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.11099999999999999, 0.135, 0.138, 0.132, 0.132, 0.138, 0.138, 0.135, 0.138, 0.135, 0.10200000000000001, 0.10800000000000001, 0.135, 0.14100000000000001, 0.138, 0.135, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.135, 0.129, 0.129, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.138, 0.15300000000000002, 0.15600000000000003, 0.22499999999999998, 0.29100000000000004, 0.339, 0.42600000000000005, 0.5309999999999999, 0.627, 0.513, 1.149, 1.077, 0.795, 0.387, 0.267, 0.21300000000000002, 0.195, 0.171, 0.165, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.132, 0.11099999999999999, 0.11399999999999999, 0.138, 0.135, 0.135, 0.11399999999999999, 0.135, 0.135, 0.132, 0.135, 0.11399999999999999, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.08700000000000001, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.11099999999999999, 0.132, 0.15600000000000003, 0.132, 0.14100000000000001, 0.15600000000000003, 0.18, 0.23399999999999999, 0.28800000000000003, 0.33, 0.393, 0.387, 0.5549999999999999, 0.81, 1.119, 0.8640000000000001, 0.396, 0.324, 0.27, 0.28800000000000003, 0.186, NaN, NaN, 0.138, 0.135, 0.138, 0.14100000000000001, 0.138, 0.135, 0.135, 0.12, 0.132, 0.129, 0.129, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.10500000000000001, 0.135, 0.132, 0.132, 0.10200000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.126, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.138, 0.14700000000000002, 0.159, 0.183, 0.22199999999999998, 0.261, 0.29400000000000004, 0.35100000000000003, 0.41700000000000004, 0.495, 0.675, 0.8550000000000001, 0.726, 0.42600000000000005, 0.44699999999999995, 0.33, 0.321, 0.31200000000000006, NaN, NaN, 0.138, 0.135, 0.135, 0.138, 0.138, 0.135, 0.138, 0.135, 0.129, 0.132, 0.11399999999999999, 0.126, 0.132, 0.138, 0.11699999999999999, 0.135, 0.081, 0.135, 0.135, 0.135, 0.138, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.132, 0.10800000000000001, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.135, 0.14700000000000002, 0.162, 0.186, 0.23099999999999998, 0.27, 0.30000000000000004, 0.28800000000000003, 0.387, 0.43799999999999994, 0.5700000000000001, 0.642, 0.726, 0.43499999999999994, 0.43200000000000005, 0.396, 0.342, 0.264, 0.321, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.126, 0.129, 0.11699999999999999, 0.135, 0.138, 0.138, 0.138, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.135, 0.11099999999999999, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.14400000000000002, 0.135, 0.14400000000000002, 0.159, 0.171, 0.21000000000000002, 0.249, 0.30000000000000004, 0.30600000000000005, 0.43799999999999994, 0.558, 0.63, 0.8699999999999999, 0.519, 0.43499999999999994, 0.366, 0.315, 0.324, NaN, NaN, 0.135, 0.135, 0.132, 0.138, 0.135, 0.138, 0.132, 0.126, 0.126, 0.132, 0.132, 0.135, 0.135, 0.132, 0.138, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.135, 0.135, 0.135, 0.10500000000000001, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.135, 0.14400000000000002, 0.15300000000000002, 0.159, 0.21899999999999997, 0.261, 0.28800000000000003, 0.255, 0.384, 0.51, 0.759, 0.759, 0.735, 0.44399999999999995, 0.366, 0.333, 0.315, 0.23399999999999999, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.138, 0.11399999999999999, 0.138, 0.138, 0.11399999999999999, 0.135, 0.129, 0.126, 0.132, 0.132, 0.14100000000000001, 0.138, 0.135, 0.138, 0.10800000000000001, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.14400000000000002, 0.165, 0.201, 0.21899999999999997, 0.273, 0.29100000000000004, 0.339, 0.387, 0.45899999999999996, 0.609, 0.741, 0.873, 0.43499999999999994, 0.35700000000000004, 0.29700000000000004, 0.30900000000000005, NaN, NaN, 0.138, 0.14100000000000001, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.138, 0.138, 0.135, 0.132, 0.129, 0.135, 0.138, 0.14100000000000001, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.10500000000000001, 0.11099999999999999, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14100000000000001, 0.15300000000000002, 0.17400000000000002, 0.20400000000000001, 0.249, 0.246, 0.276, 0.324, 0.31200000000000006, 0.396, 0.528, 0.768, 0.954, 1.332, 1.356, 0.636, 0.324, 0.28800000000000003, 0.22799999999999998, 0.246, NaN, NaN, 0.14100000000000001, 0.138, 0.135, 0.14100000000000001, 0.135, 0.135, 0.135, 0.138, 0.11399999999999999, 0.138, 0.138, 0.129, 0.14100000000000001, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.09, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.129, 0.138, 0.15000000000000002, 0.162, 0.189, 0.23399999999999999, 0.21600000000000003, 0.20700000000000002, 0.28200000000000003, 0.30600000000000005, 0.30900000000000005, 0.678, 0.8520000000000001, 1.332, 1.242, 0.9359999999999999, 0.396, 0.30600000000000005, 0.24, 0.21000000000000002, 0.21600000000000003, NaN, NaN, 0.132, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.11399999999999999, 0.129, 0.135, 0.135, 0.11099999999999999, 0.138, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.15300000000000002, 0.18, 0.237, 0.276, 0.28800000000000003, 0.327, 0.528, 0.687, 1.0050000000000001, 1.2480000000000002, 1.251, 1.287, 0.573, 0.30300000000000005, 0.261, 0.17700000000000002, 0.21899999999999997, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.138, 0.129, 0.14100000000000001, 0.135, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.14100000000000001, 0.15000000000000002, 0.171, 0.198, 0.24, 0.279, 0.318, 0.393, 0.66, 0.867, 1.0350000000000001, 1.197, 1.221, 0.891, 0.35100000000000003, 0.30900000000000005, 0.28500000000000003, 0.261, NaN, NaN, 0.138, 0.135, 0.14100000000000001, 0.138, 0.135, 0.135, 0.138, 0.135, 0.135, 0.138, 0.11099999999999999, 0.129, 0.129, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.10800000000000001, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.11399999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.10800000000000001, 0.135, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.11399999999999999, 0.14400000000000002, 0.129, 0.171, 0.189, 0.21300000000000002, 0.22499999999999998, 0.267, 0.327, 0.41700000000000004, 0.6990000000000001, 0.891, 1.131, 1.089, 0.5489999999999999, 0.42900000000000005, 0.339, 0.243, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.129, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10500000000000001, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.132, 0.132, 0.129, 0.11099999999999999, 0.138, 0.14700000000000002, 0.15300000000000002, 0.168, 0.183, 0.192, 0.22799999999999998, 0.249, 0.28500000000000003, 0.375, 0.489, 0.5820000000000001, 0.72, 0.783, 0.645, 0.489, 0.507, 0.396, 0.28800000000000003, 0.28500000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.129, 0.138, 0.132, 0.132, 0.138, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.132, 0.135, 0.12, 0.15300000000000002, 0.171, 0.189, 0.20700000000000002, 0.23099999999999998, 0.252, 0.30600000000000005, 0.366, 0.399, 0.498, 0.639, 0.756, 0.6900000000000001, 0.621, 0.399, 0.342, 0.243, 0.30300000000000005, NaN, NaN, 0.135, 0.132, 0.138, 0.138, 0.084, 0.11699999999999999, 0.135, 0.135, 0.135, 0.138, 0.10800000000000001, 0.132, 0.138, 0.132, 0.135, 0.135, 0.10800000000000001, 0.10800000000000001, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.132, 0.10500000000000001, 0.14100000000000001, 0.14700000000000002, 0.168, 0.17700000000000002, 0.17400000000000002, 0.21300000000000002, 0.237, 0.258, 0.29700000000000004, 0.40800000000000003, 0.5609999999999999, 0.666, 0.8370000000000001, 0.897, 0.8160000000000001, 0.5609999999999999, 0.43499999999999994, 0.399, 0.34500000000000003, NaN, NaN, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.135, 0.14100000000000001, 0.11399999999999999, 0.138, 0.11099999999999999, 0.135, 0.135, 0.11099999999999999, 0.129, 0.132, 0.135, 0.138, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.138, 0.129, 0.129, 0.132, 0.138, 0.14700000000000002, 0.126, 0.14400000000000002, 0.195, 0.195, 0.20400000000000001, 0.21899999999999997, 0.21000000000000002, 0.31200000000000006, 0.45899999999999996, 0.6000000000000001, 1.242, 1.362, 0.8999999999999999, 0.75, 0.43200000000000005, 0.492, 0.44399999999999995, 0.498, 0.46199999999999997, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.10800000000000001, 0.138, 0.135, 0.135, 0.11099999999999999, 0.135, 0.135, 0.132, 0.138, 0.135, 0.135, 0.132, 0.11099999999999999, 0.138, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.093, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.132, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.132, 0.138, 0.14400000000000002, 0.165, 0.17700000000000002, 0.183, 0.201, 0.23099999999999998, 0.21899999999999997, 0.46799999999999997, 0.567, 0.63, 0.7170000000000001, 0.897, 0.909, 1.059, 0.771, 0.471, 0.41700000000000004, 0.393, NaN, NaN, 0.138, 0.132, 0.138, 0.138, 0.132, 0.126, 0.126, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.138, 0.132, 0.138, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14700000000000002, 0.14400000000000002, 0.162, 0.17400000000000002, 0.189, 0.21300000000000002, 0.30000000000000004, 0.33, 0.6180000000000001, 0.639, 0.7080000000000001, 0.63, 0.5640000000000001, 1.002, 0.9510000000000001, 0.7110000000000001, 0.372, 0.28800000000000003, 0.24, 0.165, NaN, NaN, 0.135, 0.135, 0.138, 0.138, 0.138, 0.138, 0.132, 0.14100000000000001, 0.135, 0.129, 0.135, 0.14100000000000001, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.11099999999999999, 0.135, 0.11099999999999999, 0.132, 0.132, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.126, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.138, 0.14100000000000001, 0.159, 0.17700000000000002, 0.186, 0.201, 0.21300000000000002, 0.28800000000000003, 0.43200000000000005, 0.45299999999999996, 0.46199999999999997, 0.684, 0.804, 0.6060000000000001, 0.762, 0.9119999999999999, 1.1099999999999999, 0.978, 0.396, 0.324, 0.27, 0.22799999999999998, NaN, NaN, 0.138, 0.132, 0.135, 0.138, 0.11699999999999999, 0.135, 0.135, 0.135, 0.135, 0.138, 0.132, 0.132, 0.138, 0.11099999999999999, 0.135, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.10500000000000001, 0.126, 0.129, 0.129, 0.10800000000000001, 0.132, 0.135, 0.159, 0.18, 0.189, 0.17700000000000002, 0.327, 0.399, 0.44099999999999995, 0.513, 0.492, 0.519, 0.6180000000000001, 0.774, 0.996, 1.056, 0.8520000000000001, 0.498, 0.42900000000000005, 0.405, 0.327, 0.35400000000000004, 0.003, NaN, NaN, 0.138, 0.14100000000000001, 0.138, 0.132, 0.10500000000000001, 0.135, 0.123, 0.132, 0.129, 0.138, 0.14100000000000001, 0.11399999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.135, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.15300000000000002, 0.15600000000000003, 0.168, 0.168, 0.192, 0.273, 0.36, 0.46799999999999997, 0.477, 0.492, 0.474, 0.558, 0.651, 0.744, 0.75, 0.48, 0.30900000000000005, 0.381, 0.321, 0.315, 0.372, 0.43200000000000005, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.135, 0.10800000000000001, 0.135, 0.138, 0.132, 0.129, 0.129, 0.10800000000000001, 0.11399999999999999, 0.135, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.126, 0.129, 0.132, 0.135, 0.14100000000000001, 0.15000000000000002, 0.162, 0.15600000000000003, 0.168, 0.20400000000000001, 0.273, 0.336, 0.42600000000000005, 0.42900000000000005, 0.46499999999999997, 0.558, 0.627, 0.5489999999999999, 0.5760000000000001, 0.6060000000000001, 0.663, 0.513, 0.726, 0.534, 0.402, 0.384, 0.402, 0.321, 0.321, 0.387, NaN, NaN, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.129, 0.129, 0.10800000000000001, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.10500000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.10800000000000001, 0.129, 0.135, 0.129, 0.129, 0.132, 0.10800000000000001, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.159, 0.18, 0.183, 0.20700000000000002, 0.264, 0.34500000000000003, 0.41100000000000003, 0.42600000000000005, 0.5609999999999999, 0.621, 0.609, 0.5640000000000001, 0.633, 0.5549999999999999, 0.657, 0.522, 0.378, 0.369, 0.369, 0.35700000000000004, 0.30900000000000005, NaN, NaN, 0.135, 0.138, 0.138, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.126, 0.135, 0.132, 0.138, 0.135, 0.135, 0.138, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.132, 0.135, 0.14100000000000001, 0.135, 0.18, 0.17700000000000002, 0.20700000000000002, 0.28200000000000003, 0.318, 0.384, 0.471, 0.5549999999999999, 0.552, 0.41100000000000003, 0.6000000000000001, 0.522, 0.645, 0.513, 0.513, 0.372, 0.35100000000000003, 0.29700000000000004, 0.35400000000000004, 0.36, 0.279, NaN, NaN, 0.135, 0.138, 0.135, 0.132, 0.129, 0.135, 0.135, 0.132, 0.135, 0.132, 0.138, 0.11399999999999999, 0.11699999999999999, 0.135, 0.132, 0.132, 0.135, 0.135, 0.11099999999999999, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.135, 0.135, 0.138, 0.14700000000000002, 0.126, 0.168, 0.183, 0.21300000000000002, 0.29100000000000004, 0.36, 0.43499999999999994, 0.525, 0.5309999999999999, 0.54, 0.597, 0.642, 0.675, 0.579, 0.7050000000000001, 0.723, 0.5609999999999999, 0.489, 0.366, 0.36, 0.35400000000000004, 0.35400000000000004, 0.35700000000000004, 0.372, NaN, NaN, 0.138, 0.138, 0.10500000000000001, 0.135, 0.093, 0.138, 0.135, 0.135, 0.135, 0.132, 0.126, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.135, 0.138, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.129, 0.132, 0.135, 0.135, 0.138, 0.15600000000000003, 0.162, 0.18, 0.18, 0.195, 0.261, 0.35100000000000003, 0.528, 0.579, 0.669, 0.6120000000000001, 0.522, 0.627, 0.6120000000000001, 0.627, 0.474, 0.318, 0.35400000000000004, 0.35100000000000003, 0.324, 0.30900000000000005, 0.28200000000000003, NaN, NaN, 0.135, 0.126, 0.126, 0.129, 0.126, 0.129, 0.132, 0.135, 0.138, 0.135, 0.132, 0.135, 0.10200000000000001, 0.138, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.135, 0.138, 0.14100000000000001, 0.123, 0.15300000000000002, 0.168, 0.18, 0.186, 0.201, 0.22199999999999998, 0.255, 0.321, 0.375, 0.513, 0.5760000000000001, 0.6120000000000001, 0.678, 0.46799999999999997, 0.35400000000000004, 0.29100000000000004, 0.30000000000000004, 0.276, 0.237, 0.20400000000000001, 0.20400000000000001, 0.189, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.138, 0.135, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11399999999999999, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.129, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.162, 0.17400000000000002, 0.183, 0.20400000000000001, 0.22499999999999998, 0.249, 0.28200000000000003, 0.342, 0.43200000000000005, 0.46799999999999997, 0.534, 0.741, 0.492, 0.40800000000000003, 0.33, 0.342, 0.28500000000000003, 0.27, 0.252, 0.18, 0.195, 0.195, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.129, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.135, 0.129, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.11399999999999999, 0.129, 0.132, 0.132, 0.135, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.165, 0.18, 0.195, 0.22499999999999998, 0.20400000000000001, 0.279, 0.273, 0.46799999999999997, 0.43499999999999994, 0.627, 0.654, 0.78, 0.636, 0.43499999999999994, 0.399, 0.30600000000000005, 0.34500000000000003, 0.339, 0.30900000000000005, 0.23399999999999999, 0.246, NaN, NaN, 0.138, 0.126, 0.126, 0.129, 0.135, 0.132, 0.132, 0.138, 0.14100000000000001, 0.135, 0.135, 0.11399999999999999, 0.135, 0.11399999999999999, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11399999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.14100000000000001, 0.14400000000000002, 0.159, 0.171, 0.15600000000000003, 0.20400000000000001, 0.24, 0.28800000000000003, 0.34500000000000003, 0.381, 0.41400000000000003, 0.489, 0.6180000000000001, 0.687, 0.687, 0.5549999999999999, 0.34800000000000003, 0.36, 0.35100000000000003, 0.34500000000000003, 0.363, 0.35700000000000004, 0.39, 0.34500000000000003, NaN, NaN, 0.138, 0.135, 0.126, 0.126, 0.129, 0.129, 0.129, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.132, 0.09, 0.132, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.138, 0.138, 0.14700000000000002, 0.159, 0.171, 0.195, 0.20700000000000002, 0.255, 0.28200000000000003, 0.336, 0.43799999999999994, 0.495, 0.579, 0.7170000000000001, 0.675, 0.396, 0.34500000000000003, 0.372, 0.34800000000000003, 0.35100000000000003, 0.34500000000000003, 0.36, 0.342, 0.336, NaN, NaN, 0.132, 0.138, 0.135, 0.138, 0.138, 0.138, 0.138, 0.10800000000000001, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.132, 0.129, 0.11099999999999999, 0.138, 0.12, 0.165, 0.171, 0.18, 0.189, 0.198, 0.22799999999999998, 0.243, 0.273, 0.336, 0.42600000000000005, 0.5309999999999999, 0.6060000000000001, 0.7020000000000001, 0.43799999999999994, 0.34800000000000003, 0.35700000000000004, 0.35400000000000004, 0.34500000000000003, 0.336, 0.336, 0.339, NaN, NaN, 0.138, 0.138, 0.138, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.135, 0.132, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.10500000000000001, 0.132, 0.10800000000000001, 0.132, 0.135, 0.132, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.126, 0.129, 0.10800000000000001, 0.11099999999999999, 0.132, 0.14400000000000002, 0.15600000000000003, 0.165, 0.168, 0.17400000000000002, 0.15300000000000002, 0.201, 0.21899999999999997, 0.246, 0.279, 0.30900000000000005, 0.39, 0.534, 0.6120000000000001, 0.6240000000000001, 0.375, 0.342, 0.342, 0.35700000000000004, 0.339, 0.336, 0.342, NaN, NaN, 0.14100000000000001, 0.126, 0.129, 0.129, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.14100000000000001, 0.162, 0.165, 0.171, 0.192, 0.18, 0.24, 0.28500000000000003, 0.36, 0.43499999999999994, 0.579, 0.8699999999999999, 0.8490000000000001, 0.45299999999999996, 0.336, 0.33, 0.35400000000000004, 0.327, 0.27, 0.327, 0.339, NaN, NaN, 0.135, 0.132, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.129, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.09, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.14100000000000001, 0.159, 0.165, 0.183, 0.20700000000000002, 0.249, 0.267, 0.29100000000000004, 0.387, 0.45899999999999996, 0.8370000000000001, 0.8999999999999999, 0.9750000000000001, 0.768, 0.43799999999999994, 0.30900000000000005, 0.30900000000000005, 0.30600000000000005, 0.21899999999999997, 0.246, NaN, NaN, 0.135, 0.132, 0.126, 0.135, 0.135, 0.135, 0.129, 0.138, 0.138, 0.138, 0.135, 0.10800000000000001, 0.11399999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.135, 0.14100000000000001, 0.15600000000000003, 0.15600000000000003, 0.171, 0.186, 0.201, 0.186, 0.243, 0.258, 0.28200000000000003, 0.28200000000000003, 0.41700000000000004, 0.54, 0.8250000000000001, 0.7140000000000001, 0.8280000000000001, 0.678, 0.573, 0.258, 0.20700000000000002, 0.20700000000000002, 0.162, 0.192, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.138, 0.129, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.135, 0.126, 0.126, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.135, 0.14400000000000002, 0.15600000000000003, 0.15600000000000003, 0.18, 0.186, 0.20700000000000002, 0.22199999999999998, 0.249, 0.28800000000000003, 0.36, 0.44999999999999996, 0.5820000000000001, 0.879, 0.996, 0.771, 0.399, 0.29400000000000004, 0.23399999999999999, 0.168, 0.195, NaN, NaN, 0.132, 0.129, 0.10500000000000001, 0.132, 0.132, 0.132, 0.129, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.132, 0.10200000000000001, 0.132, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.129, 0.129, 0.129, 0.132, 0.135, 0.135, 0.15000000000000002, 0.14700000000000002, 0.159, 0.17400000000000002, 0.186, 0.198, 0.22199999999999998, 0.24, 0.28200000000000003, 0.384, 0.507, 0.5309999999999999, 0.9630000000000001, 1.065, 1.0050000000000001, 0.675, 0.41100000000000003, 0.35700000000000004, 0.30900000000000005, 0.261, 0.237, NaN, NaN, 0.135, 0.132, 0.135, 0.138, 0.11099999999999999, 0.138, 0.135, 0.138, 0.135, 0.135, 0.11399999999999999, 0.135, 0.11399999999999999, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.132, 0.132, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.162, 0.17700000000000002, 0.17700000000000002, 0.23099999999999998, 0.252, 0.30900000000000005, 0.31200000000000006, 0.399, 0.498, 0.732, 0.8190000000000001, 0.933, 0.8490000000000001, 0.5700000000000001, 0.474, 0.46799999999999997, 0.498, 0.489, 0.375, 0.48, NaN, NaN, 0.135, 0.135, 0.132, 0.132, 0.138, 0.138, 0.135, 0.132, 0.132, 0.132, 0.14100000000000001, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.10500000000000001, 0.09, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.138, 0.14100000000000001, 0.14700000000000002, 0.15600000000000003, 0.165, 0.192, 0.21300000000000002, 0.22199999999999998, 0.24, 0.28200000000000003, 0.33, 0.399, 0.513, 0.7170000000000001, 0.9450000000000001, 0.654, 0.621, 0.384, 0.366, 0.369, 0.336, 0.378, 0.30300000000000005, NaN, NaN, 0.135, 0.132, 0.10500000000000001, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.129, 0.11699999999999999, 0.138, 0.11399999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.132, 0.10800000000000001, 0.132, 0.14100000000000001, 0.14700000000000002, 0.162, 0.17400000000000002, 0.186, 0.201, 0.20400000000000001, 0.21300000000000002, 0.22199999999999998, 0.249, 0.29100000000000004, 0.324, 0.369, 0.46799999999999997, 0.546, 0.66, 0.8759999999999999, 0.903, 0.591, 0.30000000000000004, 0.258, 0.31200000000000006, 0.30600000000000005, 0.29400000000000004, NaN, NaN, 0.132, 0.129, 0.132, 0.132, 0.10500000000000001, 0.123, 0.126, 0.129, 0.14100000000000001, 0.138, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.10800000000000001, 0.126, 0.129, 0.10500000000000001, 0.126, 0.129, 0.135, 0.138, 0.14700000000000002, 0.14400000000000002, 0.129, 0.162, 0.183, 0.201, 0.21899999999999997, 0.246, 0.252, 0.28500000000000003, 0.34500000000000003, 0.43200000000000005, 0.522, 0.66, 0.8879999999999999, 0.642, 0.366, 0.318, 0.324, 0.318, 0.324, 0.44399999999999995, 0.402, 0.0, NaN, NaN, 0.34500000000000003, 0.333, 0.315, 0.321, 0.333, 0.327, 0.315, 0.30900000000000005, 0.31200000000000006, 0.318, 0.267, 0.318, 0.261, 0.30600000000000005, 0.30300000000000005, 0.31200000000000006, 0.30600000000000005, 0.264, 0.138, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.138, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14400000000000002, 0.15600000000000003, 0.165, 0.17700000000000002, 0.192, 0.17700000000000002, 0.201, 0.267, 0.30000000000000004, 0.36, 0.44999999999999996, 0.5489999999999999, 0.7050000000000001, 0.759, 0.43799999999999994, 0.339, 0.35100000000000003, 0.30900000000000005, 0.315, 0.30300000000000005, 0.30600000000000005, 0.30600000000000005, NaN, NaN, 0.132, 0.135, 0.11099999999999999, 0.135, 0.132, 0.135, 0.138, 0.135, 0.10800000000000001, 0.132, 0.129, 0.129, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.11099999999999999, 0.129, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.138, 0.186, 0.201, 0.22499999999999998, 0.243, 0.28500000000000003, 0.31200000000000006, 0.28500000000000003, 0.41100000000000003, 0.534, 0.879, 0.933, 0.795, 0.41100000000000003, 0.363, 0.321, 0.333, 0.29100000000000004, 0.29700000000000004, 0.273, NaN, NaN, 0.132, 0.138, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.132, 0.11399999999999999, 0.129, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.138, 0.14400000000000002, 0.15300000000000002, 0.138, 0.14700000000000002, 0.21000000000000002, 0.198, 0.261, 0.30300000000000005, 0.333, 0.363, 0.35700000000000004, 0.483, 0.567, 0.9119999999999999, 0.7050000000000001, 0.43200000000000005, 0.372, 0.35400000000000004, 0.252, 0.22799999999999998, 0.15300000000000002, 0.171, 0.159, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.10500000000000001, 0.132, 0.132, 0.08700000000000001, 0.132, 0.132, 0.135, 0.11099999999999999, 0.129, 0.132, 0.132, 0.10800000000000001, 0.126, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.15300000000000002, 0.165, 0.189, 0.22199999999999998, 0.249, 0.276, 0.30000000000000004, 0.35400000000000004, 0.327, 0.471, 0.651, 0.8400000000000001, 0.759, 0.46199999999999997, 0.363, 0.315, 0.27, 0.23399999999999999, 0.189, 0.183, 0.15600000000000003, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.138, 0.10200000000000001, 0.11099999999999999, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.135, 0.132, 0.135, 0.138, 0.11099999999999999, 0.09, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.126, 0.132, 0.129, 0.126, 0.126, 0.126, 0.132, 0.10800000000000001, 0.132, 0.138, 0.10800000000000001, 0.14700000000000002, 0.132, 0.171, 0.17700000000000002, 0.246, 0.258, 0.29100000000000004, 0.324, 0.30900000000000005, 0.42000000000000004, 0.585, 0.9870000000000001, 0.891, 0.483, 0.327, 0.30300000000000005, 0.29700000000000004, 0.261, 0.243, 0.249, 0.21899999999999997, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.10500000000000001, 0.135, 0.138, 0.135, 0.132, 0.138, 0.132, 0.11399999999999999, 0.135, 0.132, 0.11099999999999999, 0.129, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.126, 0.129, 0.10800000000000001, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.132, 0.138, 0.14700000000000002, 0.15600000000000003, 0.165, 0.171, 0.183, 0.198, 0.17700000000000002, 0.237, 0.246, 0.276, 0.342, 0.48, 0.5880000000000001, 0.8699999999999999, 1.008, 0.42000000000000004, 0.324, 0.30000000000000004, 0.28800000000000003, 0.23399999999999999, 0.27, NaN, NaN, 0.138, 0.135, 0.11099999999999999, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.10200000000000001, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.135, 0.14400000000000002, 0.15300000000000002, 0.159, 0.171, 0.186, 0.189, 0.198, 0.22799999999999998, 0.246, 0.27, 0.29400000000000004, 0.41100000000000003, 0.528, 0.573, 0.879, 0.9690000000000001, 0.42300000000000004, 0.35700000000000004, 0.34500000000000003, 0.30300000000000005, 0.279, 0.267, 0.23099999999999998, NaN, NaN, 0.138, 0.135, 0.132, 0.135, 0.135, 0.138, 0.132, 0.132, 0.11099999999999999, 0.135, 0.09, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.135, 0.11099999999999999, 0.198, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.099, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.126, 0.132, 0.132, 0.126, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.132, 0.135, 0.15000000000000002, 0.162, 0.135, 0.171, 0.195, 0.22799999999999998, 0.258, 0.28500000000000003, 0.34500000000000003, 0.46499999999999997, 0.552, 0.615, 0.8759999999999999, 0.801, 0.7050000000000001, 0.5369999999999999, 0.42300000000000004, 0.29700000000000004, 0.315, 0.273, 0.255, 0.129, NaN, NaN, 0.132, 0.138, 0.135, 0.138, 0.138, 0.135, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.138, 0.135, 0.126, 0.11399999999999999, 0.14100000000000001, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.129, 0.132, 0.138, 0.12, 0.15600000000000003, 0.159, 0.138, 0.186, 0.201, 0.237, 0.252, 0.29400000000000004, 0.378, 0.477, 0.5940000000000001, 0.8310000000000001, 0.6990000000000001, 0.792, 0.579, 0.33, 0.327, 0.29400000000000004, 0.22499999999999998, 0.264, NaN, NaN, 0.135, 0.138, 0.135, 0.135, 0.138, 0.135, 0.138, 0.132, 0.10800000000000001, 0.135, 0.135, 0.132, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.135, 0.123, 0.15300000000000002, 0.162, 0.168, 0.15600000000000003, 0.165, 0.21600000000000003, 0.23099999999999998, 0.255, 0.29700000000000004, 0.315, 0.387, 0.522, 0.753, 0.8130000000000001, 0.8759999999999999, 0.5940000000000001, 0.43200000000000005, 0.35100000000000003, 0.29700000000000004, 0.276, 0.28200000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11399999999999999, 0.11399999999999999, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.132, 0.138, 0.14700000000000002, 0.159, 0.159, 0.17400000000000002, 0.195, 0.18, 0.22199999999999998, 0.237, 0.22199999999999998, 0.28500000000000003, 0.30900000000000005, 0.363, 0.471, 0.627, 0.765, 0.909, 0.729, 0.35100000000000003, 0.243, 0.273, 0.267, 0.28500000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.10500000000000001, 0.132, 0.132, 0.126, 0.11399999999999999, 0.138, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.14400000000000002, 0.15000000000000002, 0.159, 0.183, 0.20700000000000002, 0.22199999999999998, 0.22799999999999998, 0.24, 0.255, 0.28500000000000003, 0.321, 0.372, 0.43200000000000005, 0.63, 1.032, 0.762, 0.5760000000000001, 0.35400000000000004, 0.28200000000000003, 0.246, 0.252, 0.22199999999999998, 0.21600000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.09, 0.132, 0.135, 0.132, 0.11099999999999999, 0.129, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.126, 0.129, 0.129, 0.126, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.159, 0.168, 0.171, 0.17700000000000002, 0.23399999999999999, 0.27, 0.30300000000000005, 0.375, 0.48, 0.615, 0.909, 0.783, 0.5700000000000001, 0.44399999999999995, 0.375, 0.35700000000000004, 0.30600000000000005, 0.267, 0.23399999999999999, 0.0, NaN, NaN, 0.135, 0.132, 0.135, 0.138, 0.135, 0.135, 0.138, 0.135, 0.132, 0.10800000000000001, 0.11099999999999999, 0.135, 0.11399999999999999, 0.132, 0.132, 0.126, 0.132, 0.135, 0.10800000000000001, 0.135, 0.135, 0.10500000000000001, 0.132, 0.135, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.132, 0.11099999999999999, 0.129, 0.11099999999999999, 0.10800000000000001, 0.129, 0.126, 0.129, 0.10800000000000001, 0.129, 0.126, 0.10800000000000001, 0.129, 0.126, 0.129, 0.135, 0.12, 0.15300000000000002, 0.162, 0.168, 0.14100000000000001, 0.18, 0.21000000000000002, 0.23099999999999998, 0.258, 0.31200000000000006, 0.372, 0.327, 0.525, 0.771, 0.759, 0.663, 0.489, 0.42900000000000005, 0.381, 0.321, 0.279, 0.258, 0.15600000000000003, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.132, 0.10500000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.132, 0.135, 0.129, 0.129, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.10800000000000001, 0.132, 0.10800000000000001, 0.10800000000000001, 0.132, 0.10500000000000001, 0.14400000000000002, 0.15600000000000003, 0.168, 0.18, 0.186, 0.22199999999999998, 0.252, 0.28800000000000003, 0.384, 0.402, 0.369, 0.48, 0.5489999999999999, 0.651, 0.777, 0.6960000000000001, 0.504, 0.44399999999999995, 0.41400000000000003, 0.333, 0.321, 0.30600000000000005, 0.30300000000000005, NaN, NaN, 0.135, 0.135, 0.135, 0.14100000000000001, 0.135, 0.09, 0.135, 0.138, 0.132, 0.135, 0.132, 0.132, 0.135, 0.135, 0.135, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.10800000000000001, 0.132, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.126, 0.08700000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.132, 0.10800000000000001, 0.14100000000000001, 0.15600000000000003, 0.168, 0.17700000000000002, 0.189, 0.201, 0.21600000000000003, 0.246, 0.28800000000000003, 0.264, 0.387, 0.44099999999999995, 0.492, 0.5640000000000001, 0.7050000000000001, 0.54, 0.402, 0.33, 0.29700000000000004, 0.24, 0.252, 0.31200000000000006, NaN, NaN, 0.138, 0.135, 0.132, 0.135, 0.10800000000000001, 0.135, 0.135, 0.132, 0.132, 0.135, 0.10800000000000001, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.11699999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11399999999999999, 0.10800000000000001, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.126, 0.126, 0.129, 0.129, 0.126, 0.129, 0.132, 0.14100000000000001, 0.132, 0.165, 0.18, 0.20400000000000001, 0.20700000000000002, 0.21899999999999997, 0.273, 0.336, 0.40800000000000003, 0.42300000000000004, 0.528, 0.6000000000000001, 0.675, 0.615, 0.35400000000000004, 0.369, 0.336, 0.315, 0.30000000000000004, 0.30600000000000005, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.138, 0.138, 0.093, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.126, 0.126, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.10500000000000001, 0.126, 0.126, 0.129, 0.126, 0.129, 0.11099999999999999, 0.11399999999999999, 0.14700000000000002, 0.14100000000000001, 0.17400000000000002, 0.186, 0.20700000000000002, 0.22199999999999998, 0.23399999999999999, 0.252, 0.339, 0.45599999999999996, 0.51, 0.558, 0.5549999999999999, 0.684, 0.648, 0.44099999999999995, 0.393, 0.36, 0.31200000000000006, 0.30900000000000005, 0.29100000000000004, 0.28800000000000003, NaN, NaN, 0.135, 0.135, 0.10500000000000001, 0.135, 0.132, 0.132, 0.132, 0.135, 0.11399999999999999, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.129, 0.132, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.126, 0.126, 0.10500000000000001, 0.132, 0.14700000000000002, 0.15300000000000002, 0.162, 0.17400000000000002, 0.183, 0.20400000000000001, 0.21600000000000003, 0.243, 0.267, 0.29700000000000004, 0.33, 0.519, 0.5940000000000001, 0.6990000000000001, 0.501, 0.41400000000000003, 0.35400000000000004, 0.324, 0.28200000000000003, 0.27, 0.252, 0.255, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.126, 0.129, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10500000000000001, 0.129, 0.126, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.10500000000000001, 0.138, 0.15000000000000002, 0.165, 0.17400000000000002, 0.17700000000000002, 0.159, 0.18, 0.237, 0.258, 0.261, 0.336, 0.498, 0.72, 0.6900000000000001, 0.573, 0.44099999999999995, 0.36, 0.246, 0.22799999999999998, 0.267, 0.264, 0.22199999999999998, 0.261, NaN, NaN, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.10800000000000001, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.126, 0.10800000000000001, 0.135, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.129, 0.126, 0.129, 0.129, 0.132, 0.138, 0.14700000000000002, 0.129, 0.168, 0.183, 0.201, 0.21000000000000002, 0.237, 0.27, 0.35100000000000003, 0.36, 0.501, 0.669, 0.522, 0.45299999999999996, 0.333, 0.246, 0.252, 0.22499999999999998, 0.20700000000000002, 0.17700000000000002, 0.165, 0.165, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.09, 0.132, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.08700000000000001, 0.126, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.129, 0.126, 0.129, 0.126, 0.132, 0.138, 0.15600000000000003, 0.10800000000000001, 0.17400000000000002, 0.17700000000000002, 0.195, 0.20700000000000002, 0.23399999999999999, 0.264, 0.29400000000000004, 0.333, 0.39, 0.44399999999999995, 0.663, 0.528, 0.33, 0.276, 0.21300000000000002, 0.189, 0.14400000000000002, 0.129, 0.15600000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10500000000000001, 0.129, 0.126, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.132, 0.14700000000000002, 0.15600000000000003, 0.162, 0.17400000000000002, 0.20400000000000001, 0.21600000000000003, 0.195, 0.28500000000000003, 0.34800000000000003, 0.34500000000000003, 0.486, 0.678, 0.585, 0.573, 0.35700000000000004, 0.33, 0.249, 0.23099999999999998, 0.18, 0.195, 0.183, NaN, NaN, 0.135, 0.132, 0.11399999999999999, 0.135, 0.132, 0.132, 0.138, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.126, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.129, 0.126, 0.126, 0.132, 0.14400000000000002, 0.15300000000000002, 0.162, 0.171, 0.17700000000000002, 0.195, 0.20400000000000001, 0.23099999999999998, 0.273, 0.33, 0.366, 0.45899999999999996, 0.627, 0.7080000000000001, 0.762, 0.534, 0.381, 0.28800000000000003, 0.261, 0.258, 0.255, 0.22499999999999998, 0.255, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.11399999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.126, 0.126, 0.126, 0.126, 0.10800000000000001, 0.126, 0.129, 0.132, 0.135, 0.15000000000000002, 0.15600000000000003, 0.165, 0.171, 0.192, 0.201, 0.21899999999999997, 0.258, 0.29400000000000004, 0.34500000000000003, 0.483, 0.672, 0.759, 0.654, 0.44099999999999995, 0.35100000000000003, 0.264, 0.267, 0.258, 0.255, 0.261, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.09, 0.11099999999999999, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.126, 0.123, 0.129, 0.129, 0.132, 0.14100000000000001, 0.14700000000000002, 0.138, 0.171, 0.186, 0.201, 0.20700000000000002, 0.22799999999999998, 0.24, 0.273, 0.29700000000000004, 0.372, 0.45299999999999996, 0.486, 0.639, 0.663, 0.5940000000000001, 0.42600000000000005, 0.363, 0.35100000000000003, 0.339, 0.318, 0.34800000000000003, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.126, 0.10500000000000001, 0.10800000000000001, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.10500000000000001, 0.129, 0.11399999999999999, 0.15000000000000002, 0.165, 0.17400000000000002, 0.183, 0.21300000000000002, 0.189, 0.20700000000000002, 0.30900000000000005, 0.35400000000000004, 0.42600000000000005, 0.546, 0.6000000000000001, 0.522, 0.333, 0.327, 0.31200000000000006, 0.315, 0.31200000000000006, 0.30300000000000005, 0.324, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.11399999999999999, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.126, 0.126, 0.126, 0.129, 0.126, 0.126, 0.129, 0.135, 0.11099999999999999, 0.15000000000000002, 0.165, 0.17400000000000002, 0.186, 0.165, 0.22199999999999998, 0.261, 0.29700000000000004, 0.381, 0.489, 0.603, 0.51, 0.546, 0.339, 0.44699999999999995, 0.42000000000000004, 0.504, NaN, NaN, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.10800000000000001, 0.135, 0.093, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.10500000000000001, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.10800000000000001, 0.10800000000000001, 0.126, 0.129, 0.126, 0.129, 0.10800000000000001, 0.138, 0.15000000000000002, 0.165, 0.171, 0.17400000000000002, 0.18, 0.201, 0.23399999999999999, 0.321, 0.40800000000000003, 0.44099999999999995, 0.5640000000000001, 0.7050000000000001, 0.8819999999999999, 0.5880000000000001, 0.492, 0.495, 0.78, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.135, 0.135, 0.132, 0.10200000000000001, 0.11099999999999999, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.10500000000000001, 0.129, 0.11099999999999999, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.132, 0.132, 0.135, 0.14100000000000001, 0.15000000000000002, 0.162, 0.15600000000000003, 0.171, 0.195, 0.20700000000000002, 0.21899999999999997, 0.258, 0.333, 0.321, 0.46799999999999997, 0.45599999999999996, 0.585, 0.516, 0.40800000000000003, 0.372, 0.30300000000000005, 0.315, 0.264, 0.21000000000000002, NaN, NaN, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.10800000000000001, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10500000000000001, 0.132, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.126, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10500000000000001, 0.129, 0.126, 0.08700000000000001, 0.11399999999999999, 0.129, 0.17400000000000002, 0.183, 0.192, 0.22499999999999998, 0.21000000000000002, 0.27, 0.264, 0.339, 0.522, 0.591, 0.597, 0.5309999999999999, 0.44999999999999996, 0.342, 0.333, 0.324, 0.28200000000000003, 0.29400000000000004, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.10800000000000001, 0.135, 0.132, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.138, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.10800000000000001, 0.129, 0.126, 0.129, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.135, 0.129, 0.129, 0.14400000000000002, 0.249, 0.29100000000000004, 0.28500000000000003, 0.279, 0.23399999999999999, 0.21600000000000003, 0.28200000000000003, 0.30900000000000005, 0.387, 0.36, 0.579, 0.6240000000000001, 0.498, 0.44699999999999995, 0.405, 0.336, 0.279, 0.189, NaN, NaN, 0.138, 0.135, 0.135, 0.132, 0.135, 0.10800000000000001, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.11399999999999999, 0.10800000000000001, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.132, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.126, 0.126, 0.126, 0.126, 0.129, 0.138, 0.192, 0.22199999999999998, 0.21899999999999997, 0.258, 0.28800000000000003, 0.28200000000000003, 0.29700000000000004, 0.264, 0.35100000000000003, 0.43499999999999994, 0.567, 0.645, 0.54, 0.558, 0.5369999999999999, 0.46499999999999997, 0.43499999999999994, 0.28800000000000003, NaN, NaN, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.132, 0.132, 0.14100000000000001, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.10500000000000001, 0.10800000000000001, 0.126, 0.126, 0.129, 0.10500000000000001, 0.129, 0.126, 0.126, 0.129, 0.129, 0.15300000000000002, 0.21300000000000002, 0.246, 0.21000000000000002, 0.21300000000000002, 0.252, 0.21300000000000002, 0.29100000000000004, 0.34500000000000003, 0.399, 0.41400000000000003, 0.552, 0.48, 0.333, 0.39, 0.42000000000000004, 0.44399999999999995, NaN, NaN, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.126, 0.132, 0.129, 0.10500000000000001, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.129, 0.132, 0.132, 0.135, 0.17400000000000002, 0.243, 0.201, 0.237, 0.23399999999999999, 0.279, 0.41100000000000003, 0.44999999999999996, 0.35400000000000004, 0.489, 0.489, 0.591, 0.46499999999999997, 0.43499999999999994, 0.43499999999999994, 0.46799999999999997, NaN, NaN, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.123, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.14100000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.129, 0.129, 0.129, 0.138, 0.15600000000000003, 0.237, 0.243, 0.21000000000000002, 0.22799999999999998, 0.201, 0.342, 0.591, 0.651, 0.6060000000000001, 0.44099999999999995, 0.495, 0.5369999999999999, 0.45299999999999996, 0.405, 0.318, 0.375, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.10800000000000001, 0.132, 0.135, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.10500000000000001, 0.132, 0.126, 0.126, 0.129, 0.126, 0.126, 0.10800000000000001, 0.15300000000000002, 0.135, 0.14400000000000002, 0.15300000000000002, 0.22799999999999998, 0.22799999999999998, 0.246, 0.252, 0.249, 0.264, 0.387, 0.597, 0.723, 0.8310000000000001, 0.771, 0.7050000000000001, 0.504, 0.387, 0.489, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.126, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.171, 0.129, 0.126, 0.084, 0.132, 0.126, 0.10800000000000001, 0.126, 0.126, 0.123, 0.126, 0.129, 0.10500000000000001, 0.126, 0.126, 0.11099999999999999, 0.138, 0.15000000000000002, 0.165, 0.20400000000000001, 0.255, 0.252, 0.258, 0.35100000000000003, 0.42900000000000005, 0.648, 0.762, 0.909, 0.915, 0.678, 0.507, 0.396, 0.43499999999999994, NaN, NaN, 0.138, 0.135, 0.132, 0.138, 0.10200000000000001, 0.138, 0.138, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.132, 0.129, 0.129, 0.132, 0.132, 0.135, 0.14700000000000002, 0.15300000000000002, 0.198, 0.384, 0.558, 0.522, 0.384, 0.21600000000000003, 0.195, 0.198, 0.28800000000000003, 0.41700000000000004, 0.573, 0.726, 0.645, 0.528, 0.5429999999999999, NaN, NaN, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.10800000000000001, 0.135, 0.135, 0.132, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.138, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.14100000000000001, 0.14400000000000002, 0.123, 0.14400000000000002, 0.15000000000000002, 0.165, 0.162, 0.41100000000000003, 0.684, 0.621, 0.40800000000000003, 0.399, 0.29100000000000004, 0.237, 0.22799999999999998, 0.258, 0.28500000000000003, 0.378, 0.5549999999999999, 0.75, 0.8400000000000001, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11699999999999999, 0.171, 0.30300000000000005, 0.5940000000000001, 0.6930000000000001, 0.627, 0.516, 0.46199999999999997, 0.369, 0.324, 0.276, 0.34500000000000003, 0.324, 0.585, 0.504, 0.393, NaN, NaN, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.14400000000000002, 0.132, 0.129, 0.132, 0.10500000000000001, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.14400000000000002, 0.162, 0.279, 0.378, 0.5369999999999999, 0.5700000000000001, 0.675, 0.501, 0.366, 0.30000000000000004, 0.31200000000000006, 0.36, 0.39, 0.534, 0.5429999999999999, 0.43799999999999994, 0.35100000000000003, NaN, NaN, 0.132, 0.129, 0.138, 0.132, 0.09, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.14400000000000002, 0.201, 0.22199999999999998, 0.41400000000000003, 0.642, 0.471, 0.558, 0.399, 0.28800000000000003, 0.35100000000000003, 0.41400000000000003, 0.534, 0.684, 0.771, 0.684, 0.375, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.10800000000000001, 0.138, 0.135, 0.14700000000000002, 0.183, 0.28200000000000003, 0.336, 0.678, 0.7140000000000001, 0.5940000000000001, 0.372, 0.28500000000000003, 0.45299999999999996, 0.489, 0.687, 0.897, 0.9239999999999999, 0.942, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.138, 0.11099999999999999, 0.135, 0.162, 0.22499999999999998, 0.273, 0.513, 0.654, 0.54, 0.264, 0.267, 0.381, 0.63, 0.9390000000000001, 1.119, 1.395, NaN, NaN, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11399999999999999, 0.10800000000000001, 0.132, 0.135, 0.18, 0.252, 0.31200000000000006, 0.41100000000000003, 0.633, 0.40800000000000003, 0.21000000000000002, 0.22799999999999998, 0.255, 0.558, 0.807, 1.002, 0.96, 1.0290000000000001, NaN, NaN, 0.132, 0.129, 0.129, 0.132, 0.132, 0.138, 0.132, 0.135, 0.135, 0.138, 0.192, 0.324, 0.315, 0.243, 0.5369999999999999, 0.44999999999999996, 0.138, 0.276, 0.615, 0.8939999999999999, 0.8250000000000001, 1.068, 0.942, NaN, NaN, 0.132, 0.135, 0.132, 0.135, 0.14700000000000002, 0.132, 0.129, 0.138, 0.17700000000000002, 0.249, 0.264, 0.363, 0.30000000000000004, 0.315, 0.492, 0.627, 0.471, 0.23399999999999999, 0.21300000000000002, 0.30900000000000005, 0.573, 0.774, 0.8160000000000001, 0.972, NaN, NaN, 0.138, 0.14100000000000001, 0.132, 0.14100000000000001, 0.14100000000000001, 0.138, 0.10800000000000001, 0.135, 0.135, 0.135, 0.14400000000000002, 0.15000000000000002, 0.22499999999999998, 0.33, 0.31200000000000006, 0.21600000000000003, 0.405, 0.5609999999999999, 0.636, 0.519, 0.21300000000000002, 0.267, 0.507, 0.726, 0.753, 0.8460000000000001, 0.78, NaN, NaN, 0.14700000000000002, 0.138, 0.138, 0.135, 0.138, 0.11699999999999999, 0.138, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.165, 0.276, 0.336, 0.378, 0.30900000000000005, 0.342, 0.46799999999999997, 0.5760000000000001, 0.639, 0.393, 0.318, 0.666, 0.6960000000000001, 0.723, NaN, NaN, 0.135, 0.135, 0.138, 0.138, 0.14100000000000001, 0.138, 0.135, 0.14400000000000002, 0.168, 0.162, 0.27, 0.375, 0.33, 0.255, 0.34500000000000003, 0.42300000000000004, 0.534, 0.46799999999999997, 0.237, 0.54, 0.678, 0.6900000000000001, NaN, NaN, 0.132, 0.138, 0.138, 0.138, 0.132, 0.15000000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.15600000000000003, 0.189, 0.23399999999999999, 0.315, 0.336, 0.30000000000000004, 0.279, 0.40800000000000003, 0.46199999999999997, 0.315, 0.21300000000000002, 0.327, 0.324, 0.5760000000000001, 0.591, 0.687, 0.633, NaN, NaN, 0.14400000000000002, 0.138, 0.11399999999999999, 0.138, 0.14400000000000002, 0.14400000000000002, 0.12, 0.123, 0.14700000000000002, 0.21000000000000002, 0.246, 0.30300000000000005, 0.27, 0.327, 0.483, 0.504, 0.168, 0.22799999999999998, 0.396, 0.495, 0.7080000000000001, 0.5549999999999999, NaN, NaN, 0.138, 0.135, 0.11699999999999999, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.162, 0.15000000000000002, 0.198, 0.192, 0.255, 0.36, 0.43499999999999994, 0.489, 0.387, 0.21899999999999997, 0.43799999999999994, 0.633, 0.5489999999999999, 0.633, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.123, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.186, 0.14700000000000002, 0.243, 0.315, 0.381, 0.393, 0.489, 0.483, 0.315, 0.258, 0.504, 0.657, 0.633, NaN, NaN, 0.14100000000000001, 0.138, 0.22499999999999998, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.132, 0.15300000000000002, 0.201, 0.22799999999999998, 0.267, 0.318, 0.513, 0.552, 0.30900000000000005, 0.21000000000000002, 0.31200000000000006, 0.627, 0.642, 0.5940000000000001, NaN, NaN, 0.138, 0.138, 0.123, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.15600000000000003, 0.159, 0.168, 0.201, 0.252, 0.276, 0.41400000000000003, 0.5940000000000001, 0.474, 0.20400000000000001, 0.396, 0.633, 0.609, 0.591, 0.591, 0.63, NaN, NaN, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.15300000000000002, 0.15600000000000003, 0.15300000000000002, 0.159, 0.183, 0.21600000000000003, 0.279, 0.405, 0.5369999999999999, 0.5549999999999999, 0.378, 0.18, 0.393, 0.609, 0.495, 0.552, NaN, NaN, 0.14100000000000001, 0.138, 0.14100000000000001, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.15300000000000002, 0.162, 0.138, 0.192, 0.36, 0.495, 0.5429999999999999, 0.22199999999999998, 0.246, 0.393, 0.381, 0.558, 0.42600000000000005, 0.363, 0.34500000000000003, NaN, NaN, 0.138, 0.138, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.15300000000000002, 0.14700000000000002, 0.159, 0.165, 0.168, 0.28200000000000003, 0.40800000000000003, 0.519, 0.34800000000000003, 0.342, 0.486, 0.42300000000000004, 0.477, 0.42600000000000005, 0.29700000000000004, NaN, NaN, 0.138, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.159, 0.159, 0.162, 0.171, 0.192, 0.252, 0.321, 0.46799999999999997, 0.486, 0.276, 0.44699999999999995, 0.45599999999999996, 0.522, 0.41100000000000003, 0.30900000000000005, 0.28200000000000003, NaN, NaN, 0.138, 0.14400000000000002, 0.14700000000000002, 0.15300000000000002, 0.129, 0.162, 0.15000000000000002, 0.21300000000000002, 0.21600000000000003, 0.28800000000000003, 0.44699999999999995, 0.546, 0.381, 0.273, 0.28800000000000003, 0.609, 0.43200000000000005, 0.41700000000000004, 0.318, 0.24, NaN, NaN, 0.138, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.12, 0.15000000000000002, 0.162, 0.15600000000000003, 0.183, 0.192, 0.30900000000000005, 0.522, 0.339, 0.44699999999999995, 0.507, 0.7020000000000001, 0.5700000000000001, 0.30600000000000005, 0.30600000000000005, 0.29100000000000004, NaN, NaN, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.12, 0.14700000000000002, 0.15000000000000002, 0.126, 0.165, 0.162, 0.162, 0.183, 0.21000000000000002, 0.33, 0.558, 0.663, 0.732, 0.495, 0.27, NaN, NaN, 0.138, 0.15000000000000002, 0.15600000000000003, 0.138, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.162, 0.168, 0.18, 0.186, 0.186, 0.40800000000000003, 0.498, 0.786, 0.8280000000000001, 0.384, 0.276, NaN, NaN, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.126, 0.15000000000000002, 0.15000000000000002, 0.129, 0.14400000000000002, 0.14700000000000002, 0.17400000000000002, 0.162, 0.31200000000000006, 0.41400000000000003, 0.5609999999999999, 0.8640000000000001, 0.615, 0.387, NaN, NaN, 0.138, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.126, 0.12, 0.15000000000000002, 0.135, 0.15300000000000002, 0.17400000000000002, 0.165, 0.189, 0.264, 0.405, 0.66, 0.948, 0.972, 0.678, 0.645, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.14700000000000002, 0.15300000000000002, 0.15300000000000002, 0.159, 0.159, 0.165, 0.195, 0.273, 0.519, 0.753, 0.915, 1.0530000000000002, 0.573, NaN, NaN, 0.138, 0.14400000000000002, 0.138, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.15000000000000002, 0.162, 0.138, 0.198, 0.30600000000000005, 0.35400000000000004, 0.78, 1.026, 0.8400000000000001, 0.8999999999999999, NaN, NaN, 0.14400000000000002, 0.138, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.126, 0.15000000000000002, 0.15600000000000003, 0.162, 0.138, 0.18, 0.21000000000000002, 0.372, 0.23399999999999999, 0.534, 0.684, 1.104, 0.9359999999999999, NaN, NaN, 0.14700000000000002, 0.14100000000000001, 0.15600000000000003, 0.15600000000000003, 0.171, 0.189, 0.339, 0.30300000000000005, 0.54, 0.8220000000000001, 1.1099999999999999, 0.966, 0.8580000000000001, 0.927, 0.879, 1.158, 0.891, 1.008, NaN, NaN, 0.14700000000000002, 0.15000000000000002, 0.15000000000000002, 0.159, 0.162, 0.17400000000000002, 0.252, 0.192, 0.252, 0.42600000000000005, 0.546, 0.63, 0.657, 0.726, 0.9510000000000001, 1.131, 1.104, NaN, NaN, 0.15000000000000002, 0.15300000000000002, 0.15600000000000003, 0.159, 0.15600000000000003, 0.168, 0.186, 0.24, 0.198, 0.243, 0.501, 0.573, 0.6000000000000001, 0.5609999999999999, 0.654, 0.756, 0.684, 1.014, 0.9570000000000001, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.159, 0.15000000000000002, 0.14400000000000002, 0.168, 0.135, 0.18, 0.21300000000000002, 0.43799999999999994, 0.44699999999999995, 0.657, 0.645, 0.915, 0.666, 0.8819999999999999, NaN, NaN, 0.15300000000000002, 0.15000000000000002, 0.15600000000000003, 0.15000000000000002, 0.159, 0.15600000000000003, 0.168, 0.14700000000000002, 0.14100000000000001, 0.15000000000000002, 0.171, 0.29400000000000004, 0.645, 0.948, 1.0170000000000001, 1.002, 1.044, 1.0410000000000001, 0.8520000000000001, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.15000000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.162, 0.171, 0.21300000000000002, 0.44699999999999995, 0.723, 0.933, 0.9990000000000001, 1.08, 1.113, 0.8490000000000001, 0.789, 0.8190000000000001, NaN, NaN, 0.15300000000000002, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.138, 0.15300000000000002, 0.162, 0.21300000000000002, 0.252, 0.315, 0.648, 0.8190000000000001, 0.9990000000000001, 1.089, 1.0110000000000001, 0.639, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.15000000000000002, 0.14100000000000001, 0.11699999999999999, 0.183, 0.21000000000000002, 0.21600000000000003, 0.198, 0.339, 0.573, 0.8430000000000001, 1.1219999999999999, 0.9359999999999999, 0.885, 0.885, 0.8699999999999999, NaN, NaN, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.15300000000000002, 0.165, 0.22199999999999998, 0.20400000000000001, 0.243, 0.5309999999999999, 0.798, 0.978, 0.9510000000000001, 0.8939999999999999, 0.867, 0.867, NaN, NaN, 0.14400000000000002, 0.168, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.171, 0.18, 0.18, 0.21000000000000002, 0.363, 0.615, 0.8340000000000001, 1.002, 1.026, 0.903, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.168, 0.22499999999999998, 0.35400000000000004, 0.609, 0.8759999999999999, 1.0739999999999998, 0.777, 0.774, 0.8310000000000001, 0.777, NaN, NaN, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.14100000000000001, 0.14700000000000002, 0.17700000000000002, 0.23099999999999998, 0.29400000000000004, 0.642, 0.885, 1.0739999999999998, 0.8250000000000001, 0.672, 0.6930000000000001, 0.663, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.123, 0.14100000000000001, 0.165, 0.165, 0.201, 0.30300000000000005, 0.399, 0.573, 0.9750000000000001, 1.125, 0.9990000000000001, 0.669, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.165, 0.22499999999999998, 0.35100000000000003, 0.585, 1.065, 1.0410000000000001, 0.7170000000000001, 0.6990000000000001, 0.669, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.15300000000000002, 0.135, 0.14700000000000002, 0.129, 0.21899999999999997, 0.21899999999999997, 0.381, 0.891, 0.9390000000000001, 0.7050000000000001, 0.6930000000000001, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.132, 0.138, 0.132, 0.15600000000000003, 0.168, 0.27, 0.6000000000000001, 1.068, 0.552, NaN, NaN, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.135, 0.11699999999999999, 0.14700000000000002, 0.15600000000000003, 0.336, 0.528, 0.792, 0.8879999999999999, 0.735, 0.651, 0.675, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.123, 0.135, 0.14700000000000002, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14700000000000002, 0.30600000000000005, 0.492, 0.726, 0.996, 0.786, 0.7080000000000001, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.138, 0.14400000000000002, 0.162, 0.201, 0.5369999999999999, 0.627, 0.663, 0.687, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.159, 0.17700000000000002, 0.342, 0.615, 0.885, 0.903, 0.6930000000000001, 0.585, 0.5640000000000001, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.12, 0.14700000000000002, 0.138, 0.171, 0.11399999999999999, 0.15300000000000002, 0.21000000000000002, 0.46499999999999997, 0.726, 0.9450000000000001, 0.8520000000000001, 0.681, 0.5369999999999999, 0.546, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.132, 0.14400000000000002, 0.138, 0.15000000000000002, 0.15300000000000002, 0.276, 0.6120000000000001, 0.723, 0.75, 0.489, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.14400000000000002, 0.14700000000000002, 0.123, 0.14400000000000002, 0.135, 0.14700000000000002, 0.18, 0.519, 0.63, 0.8250000000000001, 0.5760000000000001, 0.43799999999999994, 0.42300000000000004, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.11099999999999999, 0.135, 0.14700000000000002, 0.264, 0.525, 0.8190000000000001, 0.669, 0.44099999999999995, 0.375, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.138, 0.099, 0.162, 0.327, 0.5549999999999999, 0.6930000000000001, 0.366, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.138, 0.132, 0.165, 0.201, 0.40800000000000003, 0.636, 0.7140000000000001, 0.54, 0.474, 0.44099999999999995, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.135, 0.15300000000000002, 0.30000000000000004, 0.5640000000000001, 0.792, 0.669, 0.6060000000000001, 0.501, 0.45299999999999996, NaN, NaN, 0.14700000000000002, 0.14100000000000001, 0.14700000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.159, 0.30900000000000005, 0.8430000000000001, 0.6990000000000001, 0.8250000000000001, 0.507, NaN, NaN, 0.15000000000000002, 0.14700000000000002, 0.14400000000000002, 0.14700000000000002, 0.14400000000000002, 0.138, 0.15000000000000002, 0.20700000000000002, 0.525, 0.8130000000000001, 0.8580000000000001, 0.636, 0.5309999999999999, 0.42900000000000005, NaN, NaN, 0.14700000000000002, 0.14700000000000002, 0.15000000000000002, 0.14700000000000002, 0.14700000000000002, 0.138, 0.162, 0.261, 0.621, 0.741, 0.8759999999999999, 0.8160000000000001, 0.5609999999999999, 0.474, 0.42000000000000004, NaN, NaN, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.11399999999999999, 0.17400000000000002, 0.246, 0.528, 0.7050000000000001, 0.8340000000000001, 0.735, 0.5309999999999999, 0.369, NaN, NaN, 0.15000000000000002, 0.15600000000000003, 0.15000000000000002, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.43200000000000005, 0.636, 0.8699999999999999, 0.762, 0.657, 0.5640000000000001, NaN, NaN, 0.15600000000000003, 0.15300000000000002, 0.15000000000000002, 0.15300000000000002, 0.15300000000000002, 0.14100000000000001, 0.15300000000000002, 0.17400000000000002, 0.43799999999999994, 0.45599999999999996, 0.741, 0.921, 0.7020000000000001, 0.7140000000000001, 0.7110000000000001, NaN, NaN, 0.15000000000000002, 0.15000000000000002, 0.129, 0.14700000000000002, 0.14100000000000001, 0.168, 0.246, 0.579, 0.729, 0.9570000000000001, 0.8220000000000001, NaN, NaN, 0.15600000000000003, 0.162, 0.15300000000000002, 0.162, 0.132, 0.165, 0.324, 0.5309999999999999, 0.756, 0.9870000000000001, 0.8819999999999999, 0.8430000000000001, 0.8190000000000001, NaN, NaN, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.138, 0.171, 0.333, 0.5940000000000001, 0.75, 0.8999999999999999, 0.8520000000000001, 0.933, 0.8160000000000001, 0.789, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.126, 0.15300000000000002, 0.14100000000000001, 0.165, 0.28200000000000003, 0.525, 0.729, 0.8550000000000001, 0.978, 1.026, 1.05, 0.72, 0.9239999999999999, NaN, NaN, 0.17700000000000002, 0.15000000000000002, 0.15000000000000002, 0.15000000000000002, 0.29400000000000004, 0.342, 0.603, 0.774, 0.927, 1.0170000000000001, 0.8879999999999999, 0.8190000000000001, 0.8430000000000001, 0.729, NaN, NaN, 0.15600000000000003, 0.15300000000000002, 0.15300000000000002, 0.14400000000000002, 0.15000000000000002, 0.198, 0.34500000000000003, 0.54, 0.51, 0.738, 0.801, 1.002, 0.8430000000000001, 0.804, 0.867, NaN, NaN, 0.15300000000000002, 0.15300000000000002, 0.15300000000000002, 0.14700000000000002, 0.15300000000000002, 0.14100000000000001, 0.15300000000000002, 0.183, 0.333, 0.723, 0.9870000000000001, 0.8610000000000001, 0.8490000000000001, NaN, NaN, 0.15000000000000002, 0.14400000000000002, 0.15000000000000002, 0.14400000000000002, 0.14400000000000002, 0.138, 0.12, 0.15600000000000003, 0.28200000000000003, 0.9179999999999999, 0.99, 0.8939999999999999, 0.756, 0.7020000000000001, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.126, 0.14400000000000002, 0.14400000000000002, 0.18, 0.44399999999999995, 0.8939999999999999, 1.056, 0.8340000000000001, 0.744, 0.678, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.11699999999999999, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.15000000000000002, 0.186, 0.243, 0.42300000000000004, 0.615, 0.9510000000000001, 0.8610000000000001, 0.5549999999999999, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.138, 0.15000000000000002, 0.162, 0.264, 0.648, 0.762, 0.756, 0.996, 0.984, 1.056, 0.8400000000000001, 0.798, 0.8220000000000001, NaN, NaN, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.12, 0.12, 0.14400000000000002, 0.15000000000000002, 0.23399999999999999, 0.8400000000000001, 0.948, 1.1280000000000001, 1.0619999999999998, 0.9179999999999999, 0.744, 0.768, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14700000000000002, 0.14100000000000001, 0.15300000000000002, 0.14700000000000002, 0.15300000000000002, 0.17700000000000002, 0.201, 0.35700000000000004, 0.8370000000000001, 0.9810000000000001, 0.9570000000000001, 0.9810000000000001, 0.789, 0.6930000000000001, NaN, NaN, 0.138, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.138, 0.14400000000000002, 0.15000000000000002, 0.186, 0.324, 0.8460000000000001, 0.654, 0.96, 0.9239999999999999, 0.8340000000000001, 0.762, 0.744, NaN, NaN, 0.14100000000000001, 0.138, 0.138, 0.14400000000000002, 0.11099999999999999, 0.135, 0.192, 0.34500000000000003, 0.513, 0.735, 0.8699999999999999, 0.99, 1.0050000000000001, 0.8550000000000001, 0.804, 0.735, 0.7170000000000001, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.138, 0.15000000000000002, 0.14100000000000001, 0.135, 0.381, 0.5880000000000001, 0.753, 0.8640000000000001, 0.7020000000000001, 0.873, 0.6000000000000001, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.12, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.15000000000000002, 0.15300000000000002, 0.387, 0.639, 0.8939999999999999, 0.9119999999999999, 0.8999999999999999, 0.891, 0.8370000000000001, 0.8370000000000001, NaN, NaN, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14400000000000002, 0.10500000000000001, 0.138, 0.14400000000000002, 0.15300000000000002, 0.15600000000000003, 0.165, 0.165, 0.186, 0.5549999999999999, 0.792, 0.807, 0.771, 0.8190000000000001, 0.8130000000000001, NaN, NaN, 0.14100000000000001, 0.14700000000000002, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.138, 0.123, 0.138, 0.14100000000000001, 0.198, 0.30300000000000005, 0.41400000000000003, 0.7110000000000001, 0.771, 0.7170000000000001, 0.474, NaN, NaN, 0.14700000000000002, 0.14400000000000002, 0.14100000000000001, 0.138, 0.14100000000000001, 0.15000000000000002, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.165, 0.42000000000000004, 0.525, 0.741, 0.786, 0.873, 0.81, 0.72, 0.7080000000000001, 0.8340000000000001, NaN, NaN, 0.138, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.11699999999999999, 0.14400000000000002, 0.11699999999999999, 0.15300000000000002, 0.237, 0.46499999999999997, 0.603, 0.774, 0.7110000000000001, 0.807, 0.81, 0.8130000000000001, 0.7080000000000001, 0.669, 0.6900000000000001, NaN, NaN, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.15000000000000002, 0.14400000000000002, 0.14100000000000001, 0.135, 0.135, 0.14400000000000002, 0.171, 0.45599999999999996, 0.6930000000000001, 0.756, 0.807, 0.804, 0.567, 0.651, NaN, NaN, 0.135, 0.135, 0.14100000000000001, 0.14400000000000002, 0.14700000000000002, 0.15300000000000002, 0.15000000000000002, 0.162, 0.15300000000000002, 0.159, 0.165, 0.14700000000000002, 0.168, 0.22199999999999998, 0.492, 0.639, 0.768, 0.8370000000000001, 0.7020000000000001, 0.687, 0.7050000000000001, NaN, NaN, 0.15300000000000002, 0.14400000000000002, 0.14100000000000001, 0.14100000000000001, 0.14700000000000002, 0.123, 0.14700000000000002, 0.15000000000000002, 0.132, 0.15000000000000002, 0.159, 0.168, 0.21300000000000002, 0.318, 0.519, 0.684, 0.6060000000000001, 0.759, 0.669, NaN, NaN, 0.138, 0.132, 0.135, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.14700000000000002, 0.14700000000000002, 0.15300000000000002, 0.162, 0.183, 0.192, 0.198, 0.30000000000000004, 0.339, 0.28800000000000003, 0.43799999999999994, 0.44999999999999996, 0.387, 0.501, 0.558, 0.41700000000000004, 0.396, 0.399, NaN, NaN, 0.138, 0.138, 0.12, 0.138, 0.138, 0.11699999999999999, 0.15000000000000002, 0.15000000000000002, 0.162, 0.165, 0.171, 0.15300000000000002, 0.255, 0.375, 0.40800000000000003, 0.35700000000000004, 0.28200000000000003, 0.30600000000000005, 0.318, 0.42600000000000005, 0.45299999999999996, 0.363, 0.30900000000000005, NaN, NaN, 0.135, 0.132, 0.135, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.11399999999999999, 0.14700000000000002, 0.126, 0.15300000000000002, 0.162, 0.189, 0.22799999999999998, 0.31200000000000006, 0.399, 0.369, 0.23399999999999999, 0.30000000000000004, 0.40800000000000003, 0.486, 0.45899999999999996, 0.339, 0.31200000000000006, NaN, NaN, 0.132, 0.132, 0.129, 0.132, 0.14100000000000001, 0.138, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.15000000000000002, 0.15600000000000003, 0.168, 0.18, 0.21300000000000002, 0.18, 0.34500000000000003, 0.315, 0.17400000000000002, 0.267, 0.35400000000000004, 0.615, 0.75, 0.528, 0.366, NaN, NaN, 0.135, 0.135, 0.135, 0.138, 0.135, 0.11099999999999999, 0.138, 0.14400000000000002, 0.14400000000000002, 0.14400000000000002, 0.15000000000000002, 0.15000000000000002, 0.162, 0.21300000000000002, 0.23399999999999999, 0.381, 0.399, 0.20700000000000002, 0.267, 0.29400000000000004, 0.41400000000000003, 0.654, 0.5309999999999999, 0.384, 0.342, 0.33, NaN, NaN, 0.135, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.138, 0.14700000000000002, 0.15300000000000002, 0.159, 0.18, 0.198, 0.246, 0.255, 0.279, 0.35700000000000004, 0.339, 0.21899999999999997, 0.261, 0.33, 0.5700000000000001, 0.8610000000000001, 0.54, 0.33, 0.246, NaN, NaN, 0.132, 0.132, 0.129, 0.135, 0.138, 0.138, 0.138, 0.14400000000000002, 0.14700000000000002, 0.15000000000000002, 0.135, 0.18, 0.165, 0.23099999999999998, 0.36, 0.42600000000000005, 0.41400000000000003, 0.28500000000000003, 0.264, 0.35700000000000004, 0.657, 0.633, 0.759, 0.669, 0.33, NaN, NaN, 0.132, 0.132, 0.10500000000000001, 0.132, 0.135, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.14100000000000001, 0.12, 0.11399999999999999, 0.15000000000000002, 0.159, 0.195, 0.189, 0.315, 0.41100000000000003, 0.45299999999999996, 0.372, 0.34500000000000003, 0.339, 0.35100000000000003, 0.44099999999999995, 0.8430000000000001, 0.9810000000000001, 0.507, 0.42300000000000004, NaN, NaN, 0.132, 0.129, 0.135, 0.132, 0.132, 0.10800000000000001, 0.132, 0.135, 0.138, 0.138, 0.14100000000000001, 0.14400000000000002, 0.14100000000000001, 0.14400000000000002, 0.15600000000000003, 0.165, 0.198, 0.29100000000000004, 0.393, 0.44399999999999995, 0.34800000000000003, 0.31200000000000006, 0.28200000000000003, 0.31200000000000006, 0.486, 0.8759999999999999, 0.75, 0.774, 0.44399999999999995, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.135, 0.14400000000000002, 0.15300000000000002, 0.14100000000000001, 0.12, 0.14400000000000002, 0.15600000000000003, 0.20400000000000001, 0.29400000000000004, 0.34500000000000003, 0.195, 0.22199999999999998, 0.201, 0.165, 0.22499999999999998, 0.318, 0.45899999999999996, 0.762, 0.909, 0.774, 0.642, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.14700000000000002, 0.14100000000000001, 0.15300000000000002, 0.171, 0.171, 0.22199999999999998, 0.165, 0.123, 0.162, 0.14400000000000002, 0.22799999999999998, 0.339, 0.483, 0.6000000000000001, 0.777, 0.948, 0.921, 0.789, 0.789, NaN, NaN, 0.138, 0.132, 0.132, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.126, 0.10500000000000001, 0.129, 0.10200000000000001, 0.138, 0.14700000000000002, 0.162, 0.198, 0.21300000000000002, 0.33, 0.498, 0.672, 0.9179999999999999, 0.8310000000000001, 0.636, 0.729, 0.615, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.132, 0.135, 0.135, 0.135, 0.135, 0.10800000000000001, 0.132, 0.135, 0.135, 0.11099999999999999, 0.10800000000000001, 0.138, 0.135, 0.132, 0.123, 0.135, 0.138, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.135, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.129, 0.126, 0.129, 0.132, 0.135, 0.12, 0.159, 0.192, 0.22499999999999998, 0.28500000000000003, 0.336, 0.30300000000000005, 0.405, 0.525, 0.7050000000000001, 1.161, 0.663, 0.507, 0.603, NaN, NaN, 0.132, 0.132, 0.138, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.11099999999999999, 0.132, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.129, 0.126, 0.132, 0.135, 0.129, 0.132, 0.132, 0.135, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.126, 0.126, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14700000000000002, 0.171, 0.192, 0.198, 0.28500000000000003, 0.321, 0.327, 0.402, 0.363, 0.51, 0.8160000000000001, 0.903, 0.8340000000000001, 0.774, 0.8310000000000001, 0.744, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.10200000000000001, 0.135, 0.132, 0.132, 0.11399999999999999, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.126, 0.12, 0.126, 0.135, 0.132, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.135, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.132, 0.15300000000000002, 0.17700000000000002, 0.22499999999999998, 0.29700000000000004, 0.246, 0.261, 0.44099999999999995, 0.5429999999999999, 0.747, 0.8400000000000001, 0.897, 1.0619999999999998, 0.7080000000000001, 0.642, 0.735, NaN, NaN, 0.135, 0.135, 0.11399999999999999, 0.135, 0.135, 0.132, 0.138, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10500000000000001, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.18, 0.126, 0.10500000000000001, 0.126, 0.126, 0.129, 0.14400000000000002, 0.171, 0.192, 0.23399999999999999, 0.249, 0.29400000000000004, 0.44099999999999995, 0.519, 0.6240000000000001, 0.7050000000000001, 0.792, 0.6000000000000001, 0.5369999999999999, 0.35100000000000003, 0.30900000000000005, NaN, NaN, 0.135, 0.132, 0.135, 0.132, 0.11399999999999999, 0.11399999999999999, 0.135, 0.11099999999999999, 0.135, 0.11399999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.08700000000000001, 0.126, 0.129, 0.126, 0.126, 0.129, 0.10500000000000001, 0.129, 0.126, 0.129, 0.15000000000000002, 0.17400000000000002, 0.186, 0.20400000000000001, 0.21600000000000003, 0.23099999999999998, 0.23399999999999999, 0.30300000000000005, 0.45599999999999996, 0.471, 0.633, 0.7050000000000001, 0.9239999999999999, 0.777, 0.567, 0.372, 0.30300000000000005, NaN, NaN, 0.135, 0.132, 0.138, 0.138, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.10800000000000001, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.126, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.08700000000000001, 0.126, 0.126, 0.126, 0.126, 0.132, 0.129, 0.129, 0.14400000000000002, 0.15000000000000002, 0.17700000000000002, 0.195, 0.22799999999999998, 0.189, 0.189, 0.249, 0.29400000000000004, 0.34500000000000003, 0.507, 0.609, 0.765, 0.8610000000000001, 0.6930000000000001, 0.5700000000000001, 0.45299999999999996, NaN, NaN, 0.138, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.11399999999999999, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.129, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.126, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.126, 0.123, 0.126, 0.129, 0.132, 0.11399999999999999, 0.15600000000000003, 0.17700000000000002, 0.201, 0.23099999999999998, 0.24, 0.22499999999999998, 0.237, 0.318, 0.33, 0.41700000000000004, 0.567, 0.762, 1.059, 1.1400000000000001, 0.966, 0.9239999999999999, 0.726, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.10800000000000001, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.126, 0.132, 0.132, 0.129, 0.138, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.10500000000000001, 0.10500000000000001, 0.132, 0.138, 0.14400000000000002, 0.171, 0.21600000000000003, 0.23399999999999999, 0.22499999999999998, 0.22799999999999998, 0.30900000000000005, 0.29400000000000004, 0.324, 0.483, 0.66, 0.81, 0.9750000000000001, 0.867, 0.7110000000000001, 0.43499999999999994, NaN, NaN, 0.138, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.11099999999999999, 0.135, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.129, 0.129, 0.132, 0.138, 0.123, 0.165, 0.17700000000000002, 0.192, 0.23099999999999998, 0.22499999999999998, 0.23399999999999999, 0.28200000000000003, 0.393, 0.42900000000000005, 0.5940000000000001, 0.78, 1.116, 1.158, 0.744, 0.5640000000000001, 0.528, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.11399999999999999, 0.132, 0.132, 0.10500000000000001, 0.11099999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.10800000000000001, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.09, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.129, 0.132, 0.126, 0.132, 0.126, 0.129, 0.135, 0.14400000000000002, 0.171, 0.21600000000000003, 0.22199999999999998, 0.21899999999999997, 0.21300000000000002, 0.22799999999999998, 0.336, 0.381, 0.405, 0.402, 0.495, 0.534, 0.6120000000000001, 0.7170000000000001, 0.6060000000000001, 0.591, 0.567, 0.525, NaN, NaN, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.126, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.15000000000000002, 0.132, 0.129, 0.129, 0.129, 0.126, 0.10500000000000001, 0.126, 0.129, 0.126, 0.129, 0.126, 0.132, 0.129, 0.129, 0.129, 0.129, 0.11399999999999999, 0.14400000000000002, 0.162, 0.162, 0.183, 0.201, 0.22199999999999998, 0.261, 0.327, 0.381, 0.34800000000000003, 0.378, 0.43200000000000005, 0.528, 0.474, 0.5369999999999999, 0.729, 0.648, 0.615, NaN, NaN, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.11099999999999999, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.126, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.10500000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.135, 0.15000000000000002, 0.159, 0.17400000000000002, 0.186, 0.21300000000000002, 0.252, 0.31200000000000006, 0.30600000000000005, 0.29700000000000004, 0.375, 0.795, 0.9510000000000001, 1.101, 1.0230000000000001, 1.0110000000000001, 0.9690000000000001, 0.9450000000000001, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.132, 0.138, 0.132, 0.11099999999999999, 0.11099999999999999, 0.129, 0.135, 0.129, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.10500000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.138, 0.15000000000000002, 0.17700000000000002, 0.198, 0.22499999999999998, 0.264, 0.267, 0.261, 0.30600000000000005, 0.471, 0.7080000000000001, 0.7110000000000001, 0.9299999999999999, 0.9570000000000001, 0.9119999999999999, 0.639, 0.42900000000000005, NaN, NaN, 0.132, 0.138, 0.132, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.10800000000000001, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.168, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.123, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10500000000000001, 0.126, 0.126, 0.126, 0.126, 0.10800000000000001, 0.126, 0.126, 0.126, 0.129, 0.129, 0.132, 0.132, 0.14400000000000002, 0.171, 0.201, 0.23399999999999999, 0.249, 0.24, 0.21000000000000002, 0.28800000000000003, 0.30900000000000005, 0.41100000000000003, 0.5549999999999999, 0.8430000000000001, 1.083, 0.8610000000000001, 0.645, 0.43200000000000005, 0.30600000000000005, 0.249, NaN, NaN, 0.135, 0.132, 0.132, 0.132, 0.10500000000000001, 0.11099999999999999, 0.132, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.129, 0.126, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.132, 0.10800000000000001, 0.132, 0.123, 0.186, 0.22199999999999998, 0.17700000000000002, 0.21899999999999997, 0.22499999999999998, 0.237, 0.249, 0.279, 0.30000000000000004, 0.48, 0.654, 0.8610000000000001, 0.741, 0.8370000000000001, 0.672, 0.39, 0.273, NaN, NaN, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.135, 0.132, 0.11099999999999999, 0.129, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.10800000000000001, 0.132, 0.138, 0.14100000000000001, 0.15600000000000003, 0.171, 0.171, 0.171, 0.198, 0.22499999999999998, 0.22499999999999998, 0.22499999999999998, 0.246, 0.31200000000000006, 0.42600000000000005, 0.6000000000000001, 0.729, 0.8999999999999999, 0.8939999999999999, 0.879, 0.891, 0.9359999999999999, 0.756, 1.065, 1.02, NaN, NaN, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.129, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.126, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.132, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.129, 0.129, 0.132, 0.135, 0.12, 0.15300000000000002, 0.17400000000000002, 0.195, 0.22199999999999998, 0.23099999999999998, 0.24, 0.339, 0.42900000000000005, 0.5429999999999999, 0.7050000000000001, 1.221, 1.257, 1.305, 0.903, 0.789, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.10500000000000001, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.129, 0.126, 0.129, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.132, 0.135, 0.14700000000000002, 0.15600000000000003, 0.198, 0.23399999999999999, 0.237, 0.333, 0.36, 0.378, 0.48, 0.54, 0.6060000000000001, 0.63, 0.5760000000000001, 0.795, 0.897, 1.254, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.123, 0.132, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.132, 0.10800000000000001, 0.11099999999999999, 0.126, 0.129, 0.126, 0.14400000000000002, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.14100000000000001, 0.15000000000000002, 0.168, 0.198, 0.18, 0.23099999999999998, 0.255, 0.30300000000000005, 0.28800000000000003, 0.43200000000000005, 0.6240000000000001, 0.648, 1.0979999999999999, 1.1099999999999999, 1.0619999999999998, 1.158, 1.146, 0.732, 0.8939999999999999, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.10800000000000001, 0.132, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.123, 0.135, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.132, 0.129, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.126, 0.129, 0.138, 0.14700000000000002, 0.15000000000000002, 0.168, 0.186, 0.192, 0.20700000000000002, 0.261, 0.264, 0.42300000000000004, 0.603, 0.402, 0.687, 0.765, 0.8370000000000001, 0.684, 0.552, NaN, NaN, 0.132, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.099, 0.132, 0.135, 0.11099999999999999, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.126, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.135, 0.126, 0.126, 0.10800000000000001, 0.126, 0.126, 0.129, 0.126, 0.129, 0.135, 0.135, 0.135, 0.12, 0.162, 0.17700000000000002, 0.186, 0.192, 0.249, 0.30000000000000004, 0.339, 0.657, 0.5429999999999999, 0.387, 0.525, 1.0230000000000001, 0.807, 0.8250000000000001, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.129, 0.129, 0.132, 0.123, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.126, 0.126, 0.084, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.138, 0.14400000000000002, 0.159, 0.168, 0.198, 0.21300000000000002, 0.243, 0.333, 0.387, 0.777, 0.9870000000000001, 0.885, 0.8130000000000001, 0.669, 0.9990000000000001, 0.615, 0.645, NaN, NaN, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.11099999999999999, 0.132, 0.132, 0.129, 0.123, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.126, 0.126, 0.129, 0.129, 0.129, 0.132, 0.132, 0.15000000000000002, 0.15000000000000002, 0.183, 0.237, 0.252, 0.30300000000000005, 0.342, 0.34500000000000003, 0.336, 0.366, 0.46199999999999997, 0.552, 0.648, 1.368, 0.8699999999999999, 0.44399999999999995, 0.252, NaN, NaN, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.11099999999999999, 0.135, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.126, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.126, 0.10500000000000001, 0.129, 0.10500000000000001, 0.129, 0.126, 0.129, 0.129, 0.132, 0.138, 0.168, 0.189, 0.195, 0.22199999999999998, 0.21000000000000002, 0.246, 0.264, 0.28500000000000003, 0.324, 0.405, 0.41700000000000004, 0.42000000000000004, 0.663, 0.909, 0.6060000000000001, 0.34800000000000003, NaN, NaN, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.129, 0.10500000000000001, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.126, 0.126, 0.126, 0.10500000000000001, 0.126, 0.10800000000000001, 0.129, 0.129, 0.129, 0.132, 0.135, 0.135, 0.14700000000000002, 0.165, 0.162, 0.15300000000000002, 0.23399999999999999, 0.243, 0.246, 0.276, 0.36, 0.546, 0.648, 0.6060000000000001, 0.75, 1.068, 1.326, 1.1400000000000001, 0.648, NaN, NaN, 0.132, 0.135, 0.135, 0.132, 0.135, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.126, 0.135, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.126, 0.126, 0.126, 0.126, 0.10800000000000001, 0.10800000000000001, 0.129, 0.10800000000000001, 0.132, 0.132, 0.14100000000000001, 0.14400000000000002, 0.15000000000000002, 0.192, 0.237, 0.29400000000000004, 0.41700000000000004, 0.621, 0.756, 0.9810000000000001, 0.9390000000000001, 1.2240000000000002, 1.275, 1.329, 1.2240000000000002, 0.9750000000000001, 0.9450000000000001, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.135, 0.10800000000000001, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.135, 0.126, 0.129, 0.126, 0.126, 0.189, 0.129, 0.129, 0.132, 0.129, 0.129, 0.138, 0.14400000000000002, 0.14700000000000002, 0.22499999999999998, 0.243, 0.39, 0.405, 0.636, 0.8520000000000001, 0.8999999999999999, 0.9510000000000001, 0.726, 1.002, 1.0230000000000001, 1.059, 1.026, 0.8580000000000001, 0.99, NaN, NaN, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.132, 0.135, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.135, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14100000000000001, 0.15300000000000002, 0.22199999999999998, 0.27, 0.237, 0.261, 0.35700000000000004, 0.5640000000000001, 0.636, 0.678, 0.657, 0.5760000000000001, 0.723, 0.729, 0.8610000000000001, 0.6180000000000001, 0.8220000000000001, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.135, 0.135, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.132, 0.126, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.126, 0.129, 0.132, 0.138, 0.14400000000000002, 0.171, 0.249, 0.20700000000000002, 0.255, 0.33, 0.45899999999999996, 0.375, 0.5369999999999999, 0.591, 0.5549999999999999, 0.5369999999999999, 0.525, 0.867, 1.161, 1.347, 0.933, 0.8190000000000001, 0.921, NaN, NaN, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.132, 0.11099999999999999, 0.11099999999999999, 0.129, 0.132, 0.126, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.10500000000000001, 0.126, 0.10800000000000001, 0.132, 0.126, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.126, 0.129, 0.12, 0.15600000000000003, 0.198, 0.243, 0.22199999999999998, 0.30900000000000005, 0.534, 0.654, 0.42600000000000005, 0.399, 0.42600000000000005, 0.6060000000000001, 0.8340000000000001, 0.8250000000000001, 0.9870000000000001, 1.065, 0.792, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.09, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.126, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.132, 0.129, 0.14400000000000002, 0.15600000000000003, 0.22799999999999998, 0.273, 0.28500000000000003, 0.402, 0.333, 0.33, 0.375, 0.41400000000000003, 0.558, 0.765, 0.9750000000000001, 0.9059999999999999, 0.546, 0.579, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.08700000000000001, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.132, 0.123, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.132, 0.135, 0.138, 0.135, 0.192, 0.18, 0.21000000000000002, 0.237, 0.276, 0.29100000000000004, 0.30600000000000005, 0.327, 0.34800000000000003, 0.43499999999999994, 0.771, 0.8580000000000001, 0.8340000000000001, 0.741, 0.44699999999999995, 0.339, NaN, NaN, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.129, 0.11399999999999999, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.171, 0.129, 0.10800000000000001, 0.129, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.15600000000000003, 0.138, 0.11699999999999999, 0.15000000000000002, 0.186, 0.17700000000000002, 0.21000000000000002, 0.246, 0.249, 0.249, 0.249, 0.39, 0.528, 0.8220000000000001, 1.038, 0.9990000000000001, 0.66, 0.45299999999999996, 0.39, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10500000000000001, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.126, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.10800000000000001, 0.129, 0.126, 0.129, 0.132, 0.11099999999999999, 0.132, 0.138, 0.14700000000000002, 0.162, 0.189, 0.21899999999999997, 0.21899999999999997, 0.264, 0.396, 0.573, 0.9690000000000001, 0.9390000000000001, 1.125, 1.113, 1.0110000000000001, 0.8250000000000001, 0.663, NaN, NaN, 0.135, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.132, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.14100000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.135, 0.14700000000000002, 0.15000000000000002, 0.192, 0.21600000000000003, 0.22499999999999998, 0.315, 0.534, 0.636, 0.966, 1.1219999999999999, 1.161, 1.206, 1.131, 1.0619999999999998, 1.056, 0.6990000000000001, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.14100000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.129, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.10800000000000001, 0.11099999999999999, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.14100000000000001, 0.14400000000000002, 0.171, 0.195, 0.165, 0.21300000000000002, 0.35100000000000003, 0.46799999999999997, 0.546, 0.648, 0.8130000000000001, 0.9510000000000001, 1.026, 1.089, 1.095, 0.9990000000000001, 1.0110000000000001, NaN, NaN, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.132, 0.132, 0.138, 0.14400000000000002, 0.132, 0.186, 0.192, 0.29100000000000004, 0.321, 0.405, 0.516, 0.6240000000000001, 0.741, 0.804, 0.8490000000000001, 1.002, 1.092, 0.9570000000000001, 1.0290000000000001, 0.8939999999999999, 0.003, NaN, NaN, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.126, 0.129, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.138, 0.14100000000000001, 0.162, 0.189, 0.21600000000000003, 0.273, 0.30000000000000004, 0.333, 0.375, 0.44999999999999996, 0.504, 0.48, 0.498, 0.738, 1.0859999999999999, 1.0979999999999999, 0.8160000000000001, 1.194, 0.9059999999999999, 0.978, NaN, NaN, 0.132, 0.135, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.135, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.126, 0.132, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.126, 0.129, 0.10800000000000001, 0.129, 0.126, 0.129, 0.10800000000000001, 0.126, 0.10800000000000001, 0.132, 0.132, 0.135, 0.129, 0.183, 0.198, 0.243, 0.273, 0.276, 0.336, 0.363, 0.31200000000000006, 0.40800000000000003, 0.72, 1.2000000000000002, 1.314, 1.104, 0.8999999999999999, 0.75, 0.528, NaN, NaN, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.135, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.10500000000000001, 0.126, 0.132, 0.129, 0.132, 0.129, 0.10800000000000001, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.10800000000000001, 0.129, 0.129, 0.132, 0.138, 0.15300000000000002, 0.17700000000000002, 0.21899999999999997, 0.261, 0.29400000000000004, 0.28200000000000003, 0.258, 0.28500000000000003, 0.363, 0.45299999999999996, 0.44399999999999995, 0.768, 1.4220000000000002, 1.116, 1.08, 0.9179999999999999, 0.8699999999999999, 0.48, 0.34800000000000003, NaN, NaN, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.132, 0.129, 0.10500000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.11699999999999999, 0.15600000000000003, 0.14100000000000001, 0.18, 0.162, 0.198, 0.21600000000000003, 0.243, 0.28800000000000003, 0.366, 0.30600000000000005, 0.396, 0.486, 0.54, 0.948, 1.182, 0.8580000000000001, 0.75, 0.636, 0.384, 0.31200000000000006, 0.246, NaN, NaN, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.129, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.126, 0.126, 0.132, 0.129, 0.132, 0.129, 0.11099999999999999, 0.129, 0.126, 0.132, 0.10800000000000001, 0.08700000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.10800000000000001, 0.132, 0.132, 0.159, 0.165, 0.171, 0.162, 0.21600000000000003, 0.24, 0.258, 0.30600000000000005, 0.366, 0.41700000000000004, 0.471, 0.6060000000000001, 0.6240000000000001, 1.641, 0.9119999999999999, 0.8220000000000001, 0.651, 0.534, 0.471, 0.489, NaN, NaN, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.10800000000000001, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.123, 0.10500000000000001, 0.132, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.123, 0.126, 0.10500000000000001, 0.126, 0.126, 0.129, 0.132, 0.135, 0.132, 0.11699999999999999, 0.138, 0.168, 0.15300000000000002, 0.189, 0.20700000000000002, 0.23399999999999999, 0.28500000000000003, 0.342, 0.369, 0.43200000000000005, 0.522, 0.44999999999999996, 0.8759999999999999, 1.182, 1.116, 0.75, 0.738, 0.6120000000000001, 0.43799999999999994, 0.318, 0.378, NaN, NaN, 0.132, 0.129, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.129, 0.126, 0.08700000000000001, 0.129, 0.129, 0.129, 0.126, 0.126, 0.132, 0.126, 0.126, 0.126, 0.123, 0.129, 0.126, 0.126, 0.126, 0.129, 0.135, 0.14700000000000002, 0.159, 0.15300000000000002, 0.17700000000000002, 0.192, 0.201, 0.243, 0.28200000000000003, 0.33, 0.324, 0.45899999999999996, 0.5609999999999999, 0.5309999999999999, 0.46199999999999997, 0.393, 0.45599999999999996, 0.35100000000000003, 0.22499999999999998, 0.21300000000000002, 0.21300000000000002, 0.22199999999999998, 0.18, 0.165, NaN, NaN, 0.132, 0.132, 0.132, 0.138, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.132, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.123, 0.126, 0.129, 0.126, 0.126, 0.123, 0.126, 0.126, 0.132, 0.126, 0.132, 0.14100000000000001, 0.126, 0.168, 0.189, 0.21000000000000002, 0.22799999999999998, 0.249, 0.276, 0.30900000000000005, 0.342, 0.43799999999999994, 0.43499999999999994, 0.5880000000000001, 0.573, 0.726, 0.684, 0.51, 0.30600000000000005, 0.21899999999999997, 0.20700000000000002, 0.171, 0.21300000000000002, 0.11099999999999999, NaN, NaN, 0.132, 0.132, 0.14400000000000002, 0.132, 0.135, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.084, 0.126, 0.10800000000000001, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.14400000000000002, 0.15600000000000003, 0.168, 0.17700000000000002, 0.192, 0.21899999999999997, 0.24, 0.258, 0.28200000000000003, 0.33, 0.372, 0.405, 0.477, 0.495, 0.747, 0.897, 0.552, 0.28500000000000003, 0.24, 0.243, 0.279, 0.243, 0.192, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.08700000000000001, 0.129, 0.126, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.15300000000000002, 0.14700000000000002, 0.18, 0.198, 0.22199999999999998, 0.246, 0.267, 0.29400000000000004, 0.321, 0.405, 0.495, 0.5429999999999999, 0.747, 0.759, 0.327, 0.249, 0.23099999999999998, 0.22499999999999998, 0.21899999999999997, 0.22499999999999998, 0.183, 0.21899999999999997, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.123, 0.123, 0.126, 0.12, 0.126, 0.123, 0.129, 0.132, 0.14700000000000002, 0.15600000000000003, 0.18, 0.21300000000000002, 0.201, 0.28800000000000003, 0.279, 0.41400000000000003, 0.501, 0.42900000000000005, 0.7020000000000001, 0.687, 0.519, 0.369, 0.31200000000000006, 0.24, 0.24, 0.237, 0.249, 0.24, 0.24, 0.243, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.123, 0.10800000000000001, 0.10800000000000001, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.123, 0.126, 0.126, 0.10500000000000001, 0.10500000000000001, 0.126, 0.123, 0.126, 0.123, 0.126, 0.129, 0.138, 0.14400000000000002, 0.162, 0.171, 0.183, 0.195, 0.21600000000000003, 0.24, 0.264, 0.30000000000000004, 0.34800000000000003, 0.41400000000000003, 0.516, 0.666, 0.8460000000000001, 0.43200000000000005, 0.252, 0.21600000000000003, 0.252, 0.22799999999999998, 0.23399999999999999, 0.21000000000000002, 0.162, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.132, 0.10500000000000001, 0.132, 0.129, 0.129, 0.126, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.126, 0.123, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.129, 0.135, 0.138, 0.15300000000000002, 0.165, 0.11699999999999999, 0.183, 0.201, 0.23399999999999999, 0.279, 0.396, 0.495, 0.46199999999999997, 0.6120000000000001, 0.5880000000000001, 0.603, 0.255, 0.23399999999999999, 0.22499999999999998, 0.20700000000000002, 0.186, 0.18, 0.165, NaN, NaN, 0.135, 0.135, 0.132, 0.129, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.123, 0.129, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.10800000000000001, 0.126, 0.129, 0.123, 0.129, 0.126, 0.123, 0.126, 0.126, 0.132, 0.14700000000000002, 0.15300000000000002, 0.165, 0.17400000000000002, 0.189, 0.23099999999999998, 0.261, 0.327, 0.42600000000000005, 0.498, 0.546, 0.669, 0.45599999999999996, 0.276, 0.237, 0.22799999999999998, 0.22199999999999998, 0.201, 0.18, 0.171, 0.003, NaN, NaN, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.132, 0.129, 0.126, 0.129, 0.129, 0.129, 0.08700000000000001, 0.132, 0.129, 0.126, 0.126, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.123, 0.123, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.10800000000000001, 0.126, 0.135, 0.138, 0.15300000000000002, 0.168, 0.17700000000000002, 0.17700000000000002, 0.20700000000000002, 0.23399999999999999, 0.279, 0.342, 0.41100000000000003, 0.495, 0.573, 0.621, 0.45899999999999996, 0.255, 0.258, 0.249, 0.249, 0.24, 0.243, 0.24, 0.23399999999999999, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.09, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.132, 0.11099999999999999, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.135, 0.12, 0.138, 0.171, 0.15000000000000002, 0.201, 0.22199999999999998, 0.195, 0.252, 0.339, 0.42900000000000005, 0.477, 0.5609999999999999, 0.678, 0.573, 0.42300000000000004, 0.261, 0.201, 0.237, 0.246, 0.23399999999999999, 0.198, 0.23099999999999998, NaN, NaN, 0.132, 0.135, 0.10500000000000001, 0.135, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.126, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10200000000000001, 0.10500000000000001, 0.10500000000000001, 0.126, 0.126, 0.10500000000000001, 0.126, 0.129, 0.129, 0.11099999999999999, 0.14400000000000002, 0.15600000000000003, 0.168, 0.186, 0.198, 0.21300000000000002, 0.23099999999999998, 0.261, 0.321, 0.42300000000000004, 0.45599999999999996, 0.675, 0.567, 0.264, 0.249, 0.24, 0.237, 0.237, 0.23399999999999999, 0.23399999999999999, 0.23099999999999998, 0.15600000000000003, 0.237, NaN, NaN, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.10200000000000001, 0.132, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.129, 0.126, 0.10800000000000001, 0.10500000000000001, 0.126, 0.126, 0.123, 0.126, 0.123, 0.126, 0.126, 0.126, 0.132, 0.14400000000000002, 0.14100000000000001, 0.186, 0.20700000000000002, 0.22199999999999998, 0.243, 0.28500000000000003, 0.33, 0.39, 0.483, 0.507, 0.507, 0.273, 0.237, 0.237, 0.23399999999999999, 0.23399999999999999, 0.23099999999999998, 0.22799999999999998, 0.23399999999999999, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.126, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.126, 0.10500000000000001, 0.10500000000000001, 0.126, 0.123, 0.126, 0.10500000000000001, 0.126, 0.126, 0.132, 0.14400000000000002, 0.159, 0.171, 0.183, 0.198, 0.17700000000000002, 0.195, 0.258, 0.267, 0.29400000000000004, 0.33, 0.42900000000000005, 0.558, 0.687, 0.44699999999999995, 0.192, 0.22799999999999998, 0.22799999999999998, 0.22799999999999998, 0.23399999999999999, 0.23099999999999998, 0.22799999999999998, 0.22799999999999998, 0.396, NaN, NaN, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.126, 0.123, 0.11099999999999999, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.10500000000000001, 0.132, 0.126, 0.129, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.129, 0.123, 0.126, 0.126, 0.129, 0.12, 0.159, 0.159, 0.17700000000000002, 0.198, 0.23099999999999998, 0.24, 0.252, 0.29400000000000004, 0.369, 0.513, 0.5820000000000001, 0.495, 0.23399999999999999, 0.24, 0.237, 0.237, 0.24, 0.198, 0.237, 0.24, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10500000000000001, 0.132, 0.132, 0.135, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.123, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.126, 0.123, 0.123, 0.10500000000000001, 0.10500000000000001, 0.10500000000000001, 0.126, 0.126, 0.135, 0.15300000000000002, 0.168, 0.15300000000000002, 0.17700000000000002, 0.23399999999999999, 0.258, 0.28200000000000003, 0.28800000000000003, 0.387, 0.534, 0.66, 0.732, 0.45599999999999996, 0.21000000000000002, 0.21000000000000002, 0.21600000000000003, 0.17400000000000002, 0.198, 0.17700000000000002, 0.17700000000000002, 0.159, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10500000000000001, 0.129, 0.126, 0.126, 0.123, 0.126, 0.126, 0.126, 0.126, 0.132, 0.10500000000000001, 0.129, 0.138, 0.162, 0.183, 0.192, 0.18, 0.23399999999999999, 0.261, 0.31200000000000006, 0.35100000000000003, 0.42000000000000004, 0.516, 0.5940000000000001, 0.762, 0.474, 0.24, 0.23099999999999998, 0.23099999999999998, 0.21899999999999997, 0.171, 0.189, 0.18, 0.135, 0.132, 0.15600000000000003, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.132, 0.135, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.126, 0.126, 0.10800000000000001, 0.126, 0.10500000000000001, 0.126, 0.10500000000000001, 0.126, 0.123, 0.123, 0.123, 0.10500000000000001, 0.10800000000000001, 0.135, 0.14100000000000001, 0.159, 0.171, 0.186, 0.20700000000000002, 0.23399999999999999, 0.21600000000000003, 0.315, 0.375, 0.546, 0.672, 0.372, 0.246, 0.23099999999999998, 0.22499999999999998, 0.22199999999999998, 0.21300000000000002, 0.195, 0.15600000000000003, 0.171, 0.165, NaN, NaN, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.129, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.129, 0.132, 0.132, 0.129, 0.126, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.126, 0.126, 0.10500000000000001, 0.10500000000000001, 0.123, 0.123, 0.123, 0.126, 0.10500000000000001, 0.123, 0.129, 0.126, 0.10800000000000001, 0.14400000000000002, 0.129, 0.186, 0.168, 0.21600000000000003, 0.21000000000000002, 0.29100000000000004, 0.396, 0.5489999999999999, 0.558, 0.23099999999999998, 0.243, 0.243, 0.237, 0.273, 0.23399999999999999, 0.23099999999999998, 0.23099999999999998, 0.198, 0.23099999999999998, 0.23399999999999999, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.126, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.10500000000000001, 0.126, 0.126, 0.126, 0.126, 0.126, 0.10200000000000001, 0.123, 0.126, 0.10500000000000001, 0.123, 0.129, 0.129, 0.14100000000000001, 0.15000000000000002, 0.162, 0.17700000000000002, 0.183, 0.21300000000000002, 0.23099999999999998, 0.255, 0.267, 0.324, 0.471, 0.5309999999999999, 0.5700000000000001, 0.522, 0.20400000000000001, 0.246, 0.246, 0.24, 0.237, 0.249, 0.24, 0.23399999999999999, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.126, 0.123, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.12, 0.126, 0.129, 0.129, 0.126, 0.10800000000000001, 0.10500000000000001, 0.126, 0.126, 0.126, 0.123, 0.126, 0.123, 0.126, 0.126, 0.123, 0.129, 0.10800000000000001, 0.14400000000000002, 0.159, 0.14700000000000002, 0.192, 0.21600000000000003, 0.23399999999999999, 0.252, 0.321, 0.42300000000000004, 0.43499999999999994, 0.5820000000000001, 0.558, 0.36, 0.255, 0.20700000000000002, 0.249, 0.24, 0.243, 0.249, 0.252, 0.243, 0.249, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.129, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.126, 0.10800000000000001, 0.126, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.126, 0.084, 0.126, 0.126, 0.129, 0.132, 0.14400000000000002, 0.15300000000000002, 0.168, 0.186, 0.192, 0.20700000000000002, 0.22499999999999998, 0.237, 0.267, 0.339, 0.54, 0.684, 0.597, 0.246, 0.243, 0.258, 0.249, 0.246, 0.249, 0.243, 0.258, 0.246, 0.246, NaN, NaN, 0.132, 0.132, 0.10500000000000001, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.126, 0.126, 0.129, 0.129, 0.10500000000000001, 0.126, 0.129, 0.126, 0.123, 0.126, 0.084, 0.10500000000000001, 0.126, 0.10500000000000001, 0.126, 0.132, 0.135, 0.11399999999999999, 0.15300000000000002, 0.168, 0.162, 0.20700000000000002, 0.21899999999999997, 0.22799999999999998, 0.21600000000000003, 0.35400000000000004, 0.474, 0.534, 0.639, 0.5429999999999999, 0.243, 0.24, 0.237, 0.23399999999999999, 0.237, 0.23099999999999998, 0.23399999999999999, 0.23099999999999998, 0.23099999999999998, NaN, NaN, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.09, 0.129, 0.129, 0.129, 0.10800000000000001, 0.10500000000000001, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.10500000000000001, 0.10500000000000001, 0.129, 0.126, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.10200000000000001, 0.126, 0.132, 0.14700000000000002, 0.14700000000000002, 0.195, 0.171, 0.23099999999999998, 0.276, 0.336, 0.324, 0.471, 0.5309999999999999, 0.9510000000000001, 0.321, 0.23099999999999998, 0.249, 0.243, 0.237, 0.243, 0.237, 0.237, 0.201, 0.23099999999999998, 0.11099999999999999, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.10800000000000001, 0.132, 0.126, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.126, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.138, 0.123, 0.168, 0.18, 0.162, 0.20700000000000002, 0.237, 0.28500000000000003, 0.34500000000000003, 0.44699999999999995, 0.597, 0.729, 0.8190000000000001, 0.5309999999999999, 0.22499999999999998, 0.21600000000000003, 0.21300000000000002, 0.21000000000000002, 0.195, 0.183, 0.162, 0.15300000000000002, 0.14700000000000002, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.10200000000000001, 0.126, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.08700000000000001, 0.129, 0.126, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.126, 0.123, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.11099999999999999, 0.132, 0.138, 0.14700000000000002, 0.159, 0.171, 0.186, 0.195, 0.21899999999999997, 0.246, 0.30300000000000005, 0.366, 0.43799999999999994, 0.522, 0.6240000000000001, 0.9119999999999999, 0.8520000000000001, 0.366, 0.258, 0.21600000000000003, 0.20400000000000001, 0.192, 0.18, 0.162, 0.15600000000000003, 0.14400000000000002, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.129, 0.11099999999999999, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.10500000000000001, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.129, 0.126, 0.132, 0.132, 0.14100000000000001, 0.15000000000000002, 0.138, 0.17700000000000002, 0.195, 0.20400000000000001, 0.20700000000000002, 0.28800000000000003, 0.315, 0.36, 0.41100000000000003, 0.46499999999999997, 0.621, 0.897, 0.42300000000000004, 0.255, 0.23099999999999998, 0.21899999999999997, 0.195, 0.17700000000000002, 0.135, 0.15300000000000002, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.123, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.10500000000000001, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.123, 0.129, 0.126, 0.126, 0.126, 0.123, 0.126, 0.10500000000000001, 0.123, 0.126, 0.126, 0.126, 0.129, 0.132, 0.132, 0.14400000000000002, 0.159, 0.17700000000000002, 0.18, 0.192, 0.22199999999999998, 0.252, 0.30000000000000004, 0.372, 0.48, 0.8759999999999999, 0.786, 0.336, 0.29400000000000004, 0.27, 0.252, 0.21000000000000002, 0.20400000000000001, 0.24, 0.22799999999999998, 0.24, 0.22199999999999998, NaN, NaN, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.10500000000000001, 0.126, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.126, 0.10500000000000001, 0.129, 0.129, 0.129, 0.126, 0.126, 0.123, 0.126, 0.10500000000000001, 0.123, 0.126, 0.126, 0.123, 0.123, 0.126, 0.129, 0.132, 0.14700000000000002, 0.162, 0.123, 0.192, 0.22499999999999998, 0.255, 0.30300000000000005, 0.35700000000000004, 0.42600000000000005, 0.6960000000000001, 0.99, 0.42600000000000005, 0.276, 0.246, 0.23399999999999999, 0.23399999999999999, 0.23399999999999999, 0.246, 0.22799999999999998, 0.21600000000000003, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.123, 0.126, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.123, 0.126, 0.126, 0.126, 0.10500000000000001, 0.126, 0.126, 0.126, 0.08700000000000001, 0.132, 0.14100000000000001, 0.15600000000000003, 0.168, 0.165, 0.20700000000000002, 0.186, 0.23399999999999999, 0.255, 0.28200000000000003, 0.30900000000000005, 0.393, 0.5489999999999999, 0.753, 1.0110000000000001, 0.687, 0.29700000000000004, 0.29100000000000004, 0.273, 0.261, 0.243, 0.22499999999999998, 0.21899999999999997, 0.21300000000000002, 0.21899999999999997, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.123, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.10500000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.126, 0.126, 0.10500000000000001, 0.10500000000000001, 0.126, 0.126, 0.123, 0.123, 0.123, 0.10500000000000001, 0.123, 0.126, 0.126, 0.132, 0.14100000000000001, 0.129, 0.168, 0.17400000000000002, 0.189, 0.20700000000000002, 0.21600000000000003, 0.23399999999999999, 0.243, 0.279, 0.33, 0.528, 0.7020000000000001, 0.897, 0.567, 0.333, 0.29100000000000004, 0.261, 0.23399999999999999, 0.21600000000000003, 0.21300000000000002, 0.21000000000000002, 0.21000000000000002, NaN, NaN, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.126, 0.08700000000000001, 0.129, 0.126, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.123, 0.126, 0.123, 0.126, 0.126, 0.123, 0.126, 0.123, 0.10500000000000001, 0.126, 0.132, 0.11099999999999999, 0.14400000000000002, 0.165, 0.18, 0.201, 0.23099999999999998, 0.252, 0.276, 0.35100000000000003, 0.40800000000000003, 0.5429999999999999, 0.663, 0.762, 0.552, 0.318, 0.23099999999999998, 0.279, 0.28200000000000003, 0.273, 0.279, 0.22499999999999998, 0.27, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.126, 0.123, 0.135, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.126, 0.126, 0.126, 0.126, 0.126, 0.123, 0.126, 0.126, 0.123, 0.126, 0.123, 0.123, 0.126, 0.126, 0.123, 0.123, 0.123, 0.129, 0.11099999999999999, 0.132, 0.14700000000000002, 0.162, 0.18, 0.171, 0.237, 0.258, 0.24, 0.327, 0.46799999999999997, 0.666, 0.684, 0.546, 0.324, 0.28200000000000003, 0.27, 0.267, 0.255, 0.261, 0.252, 0.252, 0.249, 0.246, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.129, 0.11099999999999999, 0.132, 0.123, 0.10200000000000001, 0.135, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.132, 0.129, 0.10500000000000001, 0.126, 0.126, 0.123, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.126, 0.123, 0.126, 0.10500000000000001, 0.123, 0.123, 0.126, 0.126, 0.10500000000000001, 0.10800000000000001, 0.14100000000000001, 0.14400000000000002, 0.159, 0.17700000000000002, 0.20400000000000001, 0.183, 0.249, 0.22199999999999998, 0.321, 0.489, 0.681, 0.6930000000000001, 0.5609999999999999, 0.42600000000000005, 0.246, 0.23099999999999998, 0.21600000000000003, 0.20700000000000002, 0.189, 0.17400000000000002, 0.162, 0.15000000000000002, NaN, NaN, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.12, 0.129, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10500000000000001, 0.126, 0.126, 0.126, 0.129, 0.126, 0.126, 0.123, 0.126, 0.126, 0.126, 0.123, 0.126, 0.129, 0.099, 0.126, 0.129, 0.129, 0.11399999999999999, 0.14700000000000002, 0.15300000000000002, 0.165, 0.183, 0.21000000000000002, 0.21300000000000002, 0.246, 0.29100000000000004, 0.35100000000000003, 0.45599999999999996, 0.5489999999999999, 0.603, 0.654, 0.603, 0.396, 0.255, 0.23099999999999998, 0.22199999999999998, 0.20400000000000001, 0.195, 0.17400000000000002, 0.162, 0.159, NaN, NaN, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.123, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.10800000000000001, 0.126, 0.10500000000000001, 0.129, 0.129, 0.126, 0.126, 0.126, 0.126, 0.132, 0.10500000000000001, 0.123, 0.126, 0.099, 0.126, 0.123, 0.123, 0.126, 0.126, 0.129, 0.135, 0.11399999999999999, 0.14400000000000002, 0.15300000000000002, 0.15600000000000003, 0.186, 0.201, 0.21300000000000002, 0.21000000000000002, 0.28800000000000003, 0.35400000000000004, 0.477, 0.603, 0.6240000000000001, 0.681, 0.546, 0.30000000000000004, 0.249, 0.23099999999999998, 0.192, 0.22199999999999998, 0.21600000000000003, 0.20400000000000001, 0.201, 0.195, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.126, 0.129, 0.132, 0.10500000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.126, 0.10800000000000001, 0.126, 0.126, 0.126, 0.10200000000000001, 0.123, 0.126, 0.126, 0.126, 0.126, 0.123, 0.123, 0.126, 0.123, 0.10500000000000001, 0.129, 0.129, 0.14100000000000001, 0.15000000000000002, 0.138, 0.192, 0.20400000000000001, 0.21600000000000003, 0.24, 0.273, 0.369, 0.552, 0.639, 0.732, 0.474, 0.28500000000000003, 0.276, 0.258, 0.246, 0.243, 0.24, 0.237, 0.23099999999999998, 0.22199999999999998, 0.21600000000000003, NaN, NaN, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.126, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.11099999999999999, 0.129, 0.132, 0.10800000000000001, 0.10800000000000001, 0.10800000000000001, 0.126, 0.126, 0.126, 0.129, 0.126, 0.123, 0.123, 0.10200000000000001, 0.126, 0.123, 0.123, 0.126, 0.123, 0.126, 0.126, 0.126, 0.135, 0.15000000000000002, 0.171, 0.189, 0.198, 0.18, 0.23099999999999998, 0.276, 0.396, 0.54, 0.501, 0.42900000000000005, 0.627, 0.381, 0.17400000000000002, 0.249, 0.249, 0.237, 0.22499999999999998, 0.21899999999999997, 0.183, 0.252, NaN, NaN, 0.132, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.132, 0.126, 0.129, 0.123, 0.129, 0.135, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.126, 0.129, 0.126, 0.126, 0.126, 0.123, 0.126, 0.126, 0.123, 0.10500000000000001, 0.123, 0.12, 0.123, 0.123, 0.123, 0.126, 0.123, 0.10500000000000001, 0.132, 0.14100000000000001, 0.14400000000000002, 0.165, 0.17400000000000002, 0.192, 0.20700000000000002, 0.21899999999999997, 0.24, 0.30000000000000004, 0.396, 0.5369999999999999, 0.615, 0.519, 0.279, 0.243, 0.201, 0.23399999999999999, 0.23099999999999998, 0.23099999999999998, 0.22799999999999998, 0.22499999999999998, 0.22799999999999998, NaN, NaN, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.123, 0.123, 0.11399999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.10800000000000001, 0.126, 0.126, 0.126, 0.129, 0.10500000000000001, 0.126, 0.126, 0.126, 0.123, 0.10500000000000001, 0.123, 0.126, 0.123, 0.123, 0.126, 0.126, 0.123, 0.138, 0.129, 0.14400000000000002, 0.15000000000000002, 0.162, 0.17700000000000002, 0.198, 0.20700000000000002, 0.21899999999999997, 0.252, 0.28800000000000003, 0.35700000000000004, 0.375, 0.489, 0.552, 0.6240000000000001, 0.603, 0.321, 0.23099999999999998, 0.21600000000000003, 0.21899999999999997, 0.21899999999999997, 0.21600000000000003, 0.183, 0.18, NaN}
    DENSITY = 
      {NaN, 1026.6294, 1026.6276, 1026.6254, 1026.622, 1026.6187, 1026.6154, 1026.6104, 1026.6022, 1026.5752, 1026.5415, 1026.528, 1026.4911, 1026.4689, 1026.444, 1026.426, 1026.4192, 1026.3901, 1026.3737, 1026.3243, 1026.3032, 1026.2903, 1026.2798, 1026.2703, 1026.2546, 1026.2334, 1026.2195, 1026.201, 1026.1841, 1026.1642, 1026.1569, 1026.1499, 1026.1437, 1026.135, 1026.1274, 1026.114, 1026.0973, 1026.0695, 1026.0497, 1026.0127, 1025.973, 1025.9269, 1025.8916, 1025.8666, 1025.8531, 1025.8223, 1025.7747, 1025.7368, 1025.705, 1025.6874, 1025.6743, 1025.6543, 1025.6417, 1025.6084, 1025.5713, 1025.5461, 1025.5104, 1025.4836, 1025.4768, 1025.4689, 1025.4674, 1025.4111, 1025.4015, 1025.3627, 1025.298, 1025.2695, 1025.2338, 1025.216, 1025.2003, 1025.1775, 1025.1509, 1025.1395, 1025.1327, 1025.1274, 1025.121, 1025.1138, 1025.108, 1025.0992, 1025.0935, 1025.0869, NaN, NaN, 1026.6422, 1026.641, 1026.6381, 1026.6357, 1026.5792, 1026.5725, 1026.5492, 1026.5359, 1026.5305, 1026.5239, 1026.5168, 1026.5061, 1026.4968, 1026.4813, 1026.4617, 1026.4479, 1026.4093, 1026.3916, 1026.379, 1026.3363, 1026.3087, 1026.2946, 1026.2805, 1026.2659, 1026.2449, 1026.2346, 1026.2256, 1026.2137, 1026.2018, 1026.1606, 1026.1482, 1026.1401, 1026.1283, 1026.1198, 1026.1104, 1026.1025, 1026.0939, 1026.082, 1026.0663, 1026.0444, 1026.0332, 1026.0156, 1025.9873, 1025.9647, 1025.9202, 1025.9058, 1025.8947, 1025.8789, 1025.862, 1025.8385, 1025.8105, 1025.7828, 1025.7465, 1025.6818, 1025.6671, 1025.6201, 1025.596, 1025.5604, 1025.5306, 1025.5209, 1025.4733, 1025.4618, 1025.3854, 1025.3289, 1025.2883, 1025.2466, 1025.2308, 1025.2109, 1025.1957, 1025.1749, 1025.1677, 1025.161, 1025.1527, 1025.1466, 1025.1382, 1025.132, 1025.1266, 1025.1199, 1025.1124, 1025.1063, 1025.0935, NaN, NaN, 1026.7242, 1026.7185, 1026.7106, 1026.7035, 1026.697, 1026.6877, 1026.6776, 1026.6677, 1026.6538, 1026.6371, 1026.6084, 1026.5742, 1026.5411, 1026.5137, 1026.4684, 1026.4222, 1026.3723, 1026.3413, 1026.3143, 1026.2502, 1026.2222, 1026.1946, 1026.1682, 1026.134, 1026.1025, 1026.0507, 1026.0205, 1025.9777, 1025.9155, 1025.871, 1025.817, 1025.7198, 1025.6455, 1025.5824, 1025.494, 1025.3955, 1025.3192, 1025.2341, 1025.2125, 1025.1986, 1025.186, 1025.1737, 1025.1594, 1025.1454, 1025.1273, 1025.1149, 1025.0999, NaN, NaN, 1026.8013, 1026.7883, 1026.7742, 1026.7473, 1026.7245, 1026.715, 1026.705, 1026.6938, 1026.681, 1026.6664, 1026.6548, 1026.6432, 1026.628, 1026.6134, 1026.59, 1026.574, 1026.5463, 1026.5227, 1026.5034, 1026.413, 1026.344, 1026.3204, 1026.254, 1026.2184, 1026.1853, 1026.1573, 1026.1377, 1026.1097, 1026.0602, 1026.0183, 1025.9534, 1025.9169, 1025.8739, 1025.8303, 1025.7312, 1025.66, 1025.5898, 1025.4866, 1025.4144, 1025.3455, 1025.2314, 1025.2148, 1025.2002, 1025.1868, 1025.1661, 1025.1335, 1025.0831, 1025.0261, 1025.0029, 1024.9772, NaN, NaN, 1026.8262, 1026.8201, 1026.8033, 1026.7843, 1026.7684, 1026.7534, 1026.7289, 1026.7163, 1026.7018, 1026.6863, 1026.6731, 1026.6592, 1026.6437, 1026.6228, 1026.592, 1026.5117, 1026.4633, 1026.4227, 1026.3788, 1026.363, 1026.3483, 1026.327, 1026.2776, 1026.2495, 1026.2213, 1026.196, 1026.1666, 1026.1326, 1026.1017, 1026.0311, 1025.9795, 1025.9432, 1025.8981, 1025.8528, 1025.8059, 1025.733, 1025.6364, 1025.546, 1025.4551, 1025.3977, 1025.3499, 1025.2499, 1025.2277, 1025.2109, 1025.1998, 1025.1792, 1025.1566, 1025.1332, 1025.0936, 1025.0089, 1024.987, 1024.9591, NaN, NaN, 1026.8627, 1026.8475, 1026.8329, 1026.8137, 1026.7893, 1026.7755, 1026.7645, 1026.7545, 1026.7421, 1026.73, 1026.7195, 1026.7076, 1026.6953, 1026.6753, 1026.6293, 1026.605, 1026.5574, 1026.534, 1026.5092, 1026.4883, 1026.4581, 1026.404, 1026.3593, 1026.3333, 1026.3165, 1026.2869, 1026.2406, 1026.2042, 1026.1764, 1026.1251, 1026.0458, 1026.0095, 1025.9912, 1025.9757, 1025.949, 1025.8851, 1025.8362, 1025.7651, 1025.6981, 1025.6165, 1025.5204, 1025.4729, 1025.4362, 1025.4037, 1025.3408, 1025.2361, 1025.205, 1025.1888, 1025.1736, 1025.1428, 1025.103, 1025.0039, 1024.9539, 1024.9368, 1024.9218, 1024.906, NaN, NaN, 1026.8622, 1026.8488, 1026.8427, 1026.8276, 1026.8175, 1026.8079, 1026.797, 1026.7809, 1026.7504, 1026.7233, 1026.7029, 1026.6765, 1026.6611, 1026.6432, 1026.6213, 1026.6062, 1026.5762, 1026.5568, 1026.5317, 1026.5051, 1026.4719, 1026.4191, 1026.384, 1026.3511, 1026.3032, 1026.2662, 1026.2404, 1026.2153, 1026.1669, 1026.1246, 1026.0917, 1026.0499, 1025.9906, 1025.9749, 1025.9634, 1025.9547, 1025.9268, 1025.8468, 1025.7975, 1025.7549, 1025.6774, 1025.6088, 1025.5468, 1025.4945, 1025.443, 1025.3955, 1025.3514, 1025.2723, 1025.195, 1025.1687, 1025.1364, 1025.0712, 1025.0098, 1024.9398, 1024.925, 1024.9061, NaN, NaN, 1026.8943, 1026.8728, 1026.8616, 1026.8507, 1026.8387, 1026.8234, 1026.8065, 1026.7881, 1026.7588, 1026.7289, 1026.7069, 1026.6761, 1026.6309, 1026.5828, 1026.538, 1026.4926, 1026.4666, 1026.4515, 1026.4309, 1026.4083, 1026.3601, 1026.3243, 1026.3102, 1026.2888, 1026.2579, 1026.2333, 1026.2085, 1026.1864, 1026.1439, 1026.1229, 1026.1006, 1026.0049, 1025.9158, 1025.8693, 1025.8142, 1025.7789, 1025.7467, 1025.7162, 1025.6353, 1025.58, 1025.5386, 1025.4426, 1025.4081, 1025.3833, 1025.3503, 1025.2782, 1025.244, 1025.1885, 1025.1373, 1025.0922, 1025.0238, 1024.9565, 1024.9414, 1024.9254, 1024.8969, 1024.8657, NaN, NaN, 1026.9231, 1026.9176, 1026.904, 1026.8903, 1026.8763, 1026.8604, 1026.8463, 1026.8356, 1026.8135, 1026.7928, 1026.7595, 1026.7308, 1026.6945, 1026.6681, 1026.6298, 1026.6005, 1026.5771, 1026.537, 1026.5028, 1026.4684, 1026.4484, 1026.4355, 1026.4155, 1026.3896, 1026.3463, 1026.3297, 1026.312, 1026.2698, 1026.2385, 1026.2205, 1026.1849, 1026.1621, 1026.1295, 1026.0437, 1025.953, 1025.8951, 1025.8507, 1025.8104, 1025.7505, 1025.6671, 1025.6061, 1025.5406, 1025.472, 1025.3916, 1025.3672, 1025.3226, 1025.2367, 1025.1874, 1025.1542, 1025.1089, 1025.0895, 1025.0746, 1024.9775, 1024.953, 1024.9415, 1024.9331, 1024.9031, 1024.8845, 1024.8706, 1024.8119, NaN, NaN, 1026.9628, 1026.956, 1026.9506, 1026.9375, 1026.9274, 1026.9153, 1026.9048, 1026.8914, 1026.8728, 1026.8431, 1026.826, 1026.7982, 1026.7632, 1026.7411, 1026.7073, 1026.6779, 1026.6348, 1026.606, 1026.5835, 1026.5646, 1026.5411, 1026.5054, 1026.4702, 1026.4479, 1026.4233, 1026.3744, 1026.325, 1026.2853, 1026.2538, 1026.2216, 1026.1915, 1026.1636, 1026.0382, 1025.9478, 1025.8975, 1025.8757, 1025.8508, 1025.8157, 1025.7922, 1025.7642, 1025.7358, 1025.7173, 1025.6819, 1025.6086, 1025.5715, 1025.5433, 1025.4733, 1025.4447, 1025.4028, 1025.3329, 1025.3064, 1025.2583, 1025.1366, 1025.0316, 1024.9492, 1024.9241, 1024.9055, 1024.8679, 1024.8235, 1024.7802, 1024.754, 1024.7319, NaN, NaN, 1026.9921, 1026.986, 1026.975, 1026.966, 1026.9565, 1026.9448, 1026.9343, 1026.9235, 1026.9065, 1026.8856, 1026.865, 1026.8469, 1026.8251, 1026.8041, 1026.7797, 1026.7528, 1026.7249, 1026.6912, 1026.6681, 1026.6489, 1026.627, 1026.6075, 1026.575, 1026.534, 1026.4948, 1026.4609, 1026.4061, 1026.3868, 1026.3679, 1026.3019, 1026.2628, 1026.2245, 1026.1886, 1026.1538, 1026.106, 1025.9862, 1025.947, 1025.9222, 1025.9086, 1025.8884, 1025.7866, 1025.7173, 1025.6921, 1025.6724, 1025.6295, 1025.563, 1025.509, 1025.449, 1025.3538, 1025.2953, 1025.2399, 1025.1733, 1025.102, 1024.9987, 1024.9636, 1024.9156, 1024.8408, 1024.8086, 1024.7777, 1024.7374, 1024.7047, 1024.6747, NaN, NaN, 1027.0419, 1027.0343, 1027.0287, 1027.0189, 1027.01, 1027.0, 1026.9901, 1026.9791, 1026.9652, 1026.947, 1026.9321, 1026.9187, 1026.8949, 1026.8694, 1026.8433, 1026.8273, 1026.8108, 1026.7853, 1026.7532, 1026.7318, 1026.7025, 1026.6792, 1026.6614, 1026.6365, 1026.6141, 1026.5789, 1026.5359, 1026.493, 1026.4552, 1026.4191, 1026.3849, 1026.344, 1026.3229, 1026.3008, 1026.2578, 1026.2207, 1026.1974, 1026.1678, 1026.1077, 1026.0625, 1025.9801, 1025.9564, 1025.9326, 1025.9077, 1025.8748, 1025.8232, 1025.7081, 1025.6228, 1025.5745, 1025.5509, 1025.4943, 1025.4266, 1025.305, 1025.2526, 1025.2174, 1025.1764, 1025.1149, 1025.0687, 1025.034, 1024.9861, 1024.9475, 1024.8835, 1024.7894, 1024.7513, 1024.7354, 1024.7163, NaN, NaN, 1027.1343, 1027.1208, 1027.1056, 1027.0874, 1027.0585, 1027.0258, 1026.996, 1026.967, 1026.9376, 1026.9064, 1026.8677, 1026.8358, 1026.7924, 1026.7678, 1026.7166, 1026.676, 1026.6127, 1026.5349, 1026.4625, 1026.3829, 1026.3156, 1026.2229, 1026.1024, 1026.0297, 1025.9706, 1025.9169, 1025.749, 1025.5907, 1025.5242, 1025.4719, 1025.3422, 1025.2609, 1025.1477, 1025.076, 1025.0298, 1024.889, 1024.8123, 1024.7715, 1024.7565, NaN, NaN, 1027.3405, 1027.3079, 1027.2638, 1027.2166, 1027.1625, 1027.1235, 1027.0905, 1027.0543, 1027.0193, 1026.9825, 1026.9463, 1026.9099, 1026.8723, 1026.8235, 1026.7832, 1026.7391, 1026.6799, 1026.6052, 1026.5073, 1026.4393, 1026.3734, 1026.313, 1026.2338, 1026.183, 1026.1132, 1026.0566, 1025.9917, 1025.9395, 1025.8651, 1025.6843, 1025.5891, 1025.4656, 1025.371, 1025.2515, 1025.1652, 1025.1238, 1025.0452, 1024.9608, 1024.8752, 1024.8188, NaN, NaN, 1027.5461, 1027.528, 1027.4745, 1027.417, 1027.3682, 1027.3318, 1027.2781, 1027.2264, 1027.1855, 1027.1362, 1027.1017, 1027.069, 1027.032, 1026.9966, 1026.9639, 1026.9127, 1026.8613, 1026.8007, 1026.7473, 1026.684, 1026.6213, 1026.542, 1026.4875, 1026.4454, 1026.3976, 1026.3422, 1026.2848, 1026.1948, 1026.1249, 1026.068, 1026.0127, 1025.9408, 1025.9036, 1025.8519, 1025.7661, 1025.6274, 1025.4706, 1025.3635, 1025.2933, 1025.2169, 1025.1472, 1025.1143, 1025.0287, 1024.893, 1024.7969, NaN, NaN, 1027.7437, 1027.7295, 1027.7122, 1027.6946, 1027.6713, 1027.6511, 1027.6301, 1027.6072, 1027.5748, 1027.5114, 1027.4678, 1027.4226, 1027.3569, 1027.2938, 1027.2543, 1027.2062, 1027.1534, 1027.1111, 1027.0769, 1027.0253, 1026.9777, 1026.9424, 1026.9164, 1026.8911, 1026.8623, 1026.827, 1026.8002, 1026.7477, 1026.6863, 1026.6564, 1026.5917, 1026.5189, 1026.4899, 1026.4606, 1026.4022, 1026.349, 1026.2677, 1026.1583, 1026.0391, 1025.9215, 1025.8773, 1025.712, 1025.5898, 1025.4965, 1025.4249, 1025.3508, 1025.2883, 1025.1752, 1025.0906, 1025.046, 1025.0076, 1024.9753, 1024.9159, 1024.8655, NaN, NaN, 1027.8553, 1027.8363, 1027.8118, 1027.7822, 1027.7401, 1027.6952, 1027.6448, 1027.6018, 1027.5587, 1027.5216, 1027.4778, 1027.4288, 1027.3721, 1027.3307, 1027.3004, 1027.2626, 1027.2239, 1027.1631, 1027.124, 1027.0863, 1027.0541, 1027.0197, 1026.963, 1026.9102, 1026.8743, 1026.8165, 1026.7524, 1026.6875, 1026.6359, 1026.574, 1026.507, 1026.4297, 1026.351, 1026.3123, 1026.256, 1026.2013, 1026.1631, 1026.02, 1025.9487, 1025.8959, 1025.8177, 1025.6726, 1025.5497, 1025.4631, 1025.3019, 1025.2429, 1025.1345, 1025.0493, 1024.9908, 1024.9318, 1024.8503, 1024.7458, NaN, NaN, 1027.9778, 1027.9635, 1027.9451, 1027.9196, 1027.889, 1027.8625, 1027.8263, 1027.7947, 1027.7576, 1027.7122, 1027.6635, 1027.6373, 1027.6082, 1027.5737, 1027.5321, 1027.4921, 1027.4519, 1027.4182, 1027.3683, 1027.3346, 1027.2781, 1027.2301, 1027.1816, 1027.1313, 1027.0967, 1027.0582, 1027.0105, 1026.9679, 1026.9153, 1026.863, 1026.8353, 1026.8004, 1026.7463, 1026.6731, 1026.5985, 1026.5339, 1026.465, 1026.4126, 1026.3694, 1026.3279, 1026.2917, 1026.2422, 1026.1942, 1026.156, 1026.1083, 1026.0599, 1025.9554, 1025.8193, 1025.7086, 1025.5956, 1025.51, 1025.4435, 1025.3114, 1025.197, 1024.9912, 1024.9541, 1024.911, 1024.8833, 1024.8279, 1024.7686, 1024.6803, NaN, NaN, 1028.2102, 1028.197, 1028.1766, 1028.1464, 1028.1075, 1028.0701, 1028.0392, 1028.0148, 1027.9895, 1027.9612, 1027.9338, 1027.9058, 1027.8727, 1027.8376, 1027.8064, 1027.7771, 1027.7476, 1027.705, 1027.6763, 1027.6514, 1027.6084, 1027.5725, 1027.5208, 1027.4866, 1027.4625, 1027.4362, 1027.392, 1027.3529, 1027.3204, 1027.2861, 1027.2416, 1027.1998, 1027.1477, 1027.0984, 1027.0618, 1027.0094, 1026.9463, 1026.9004, 1026.8557, 1026.8279, 1026.7731, 1026.7122, 1026.6622, 1026.6079, 1026.5459, 1026.4562, 1026.3722, 1026.346, 1026.313, 1026.2681, 1026.2343, 1026.2056, 1026.162, 1026.1023, 1026.0477, 1025.9553, 1025.8617, 1025.7384, 1025.6752, 1025.5497, 1025.3888, 1025.318, 1025.2234, 1025.1295, 1025.0028, 1024.9152, 1024.8772, 1024.841, 1024.7737, 1024.6921, 1024.6417, NaN, NaN, 1028.5712, 1028.55, 1028.5186, 1028.4951, 1028.4717, 1028.4476, 1028.4169, 1028.3877, 1028.3541, 1028.3141, 1028.2733, 1028.2334, 1028.1993, 1028.1699, 1028.1357, 1028.1031, 1028.0728, 1028.0319, 1027.9852, 1027.9539, 1027.9119, 1027.8794, 1027.8472, 1027.8126, 1027.7753, 1027.7452, 1027.7096, 1027.6809, 1027.6442, 1027.5945, 1027.549, 1027.5013, 1027.4674, 1027.43, 1027.3884, 1027.3495, 1027.3165, 1027.2742, 1027.2229, 1027.1787, 1027.1282, 1027.0679, 1027.0269, 1026.9613, 1026.8806, 1026.8009, 1026.7664, 1026.7249, 1026.6633, 1026.6075, 1026.5509, 1026.5061, 1026.4508, 1026.3965, 1026.3618, 1026.3013, 1026.2506, 1026.1486, 1026.0742, 1025.9994, 1025.9235, 1025.8087, 1025.7377, 1025.6423, 1025.5264, 1025.4185, 1025.2633, 1025.207, 1025.1067, 1024.9402, 1024.8683, 1024.8453, 1024.7777, 1024.7207, 1024.6794, 1024.6215, 1024.5614, NaN, NaN, 1028.6406, 1028.6276, 1028.5845, 1028.5552, 1028.5138, 1028.478, 1028.4385, 1028.3936, 1028.3606, 1028.3265, 1028.2828, 1028.2402, 1028.2075, 1028.1746, 1028.1427, 1028.1096, 1028.0754, 1028.046, 1027.9976, 1027.9672, 1027.925, 1027.885, 1027.8524, 1027.8188, 1027.7882, 1027.7482, 1027.7087, 1027.6711, 1027.6345, 1027.598, 1027.5505, 1027.5173, 1027.4868, 1027.4569, 1027.4281, 1027.3944, 1027.3638, 1027.3291, 1027.2952, 1027.2612, 1027.2249, 1027.191, 1027.1466, 1027.1007, 1027.0465, 1026.973, 1026.9357, 1026.8914, 1026.8411, 1026.7808, 1026.73, 1026.6425, 1026.6036, 1026.5538, 1026.503, 1026.4233, 1026.3652, 1026.3281, 1026.2748, 1026.2278, 1026.1827, 1026.1228, 1026.0753, 1025.952, 1025.8921, 1025.7848, 1025.7114, 1025.5991, 1025.5283, 1025.4332, 1025.2854, 1025.1278, 1025.0759, 1024.9636, 1024.8527, 1024.8308, 1024.8005, 1024.7463, 1024.67, 1024.594, 1024.567, NaN, NaN, 1028.5557, 1028.5417, 1028.5209, 1028.5029, 1028.4641, 1028.4318, 1028.3978, 1028.3633, 1028.3317, 1028.2965, 1028.2657, 1028.221, 1028.1884, 1028.1589, 1028.1161, 1028.0771, 1028.0414, 1028.0111, 1027.9834, 1027.9575, 1027.9286, 1027.895, 1027.8584, 1027.8263, 1027.794, 1027.7659, 1027.7347, 1027.7009, 1027.6697, 1027.6361, 1027.6024, 1027.5724, 1027.5348, 1027.5029, 1027.4667, 1027.4355, 1027.3918, 1027.3605, 1027.3275, 1027.2882, 1027.2495, 1027.1927, 1027.153, 1027.1108, 1027.0822, 1027.0435, 1026.9819, 1026.9365, 1026.8956, 1026.8511, 1026.7908, 1026.7362, 1026.6876, 1026.6167, 1026.556, 1026.47, 1026.4069, 1026.3663, 1026.303, 1026.2072, 1026.1383, 1026.0806, 1026.0114, 1025.9398, 1025.8394, 1025.7588, 1025.6849, 1025.5935, 1025.4988, 1025.3541, 1025.2103, 1024.9642, 1024.9116, 1024.8578, 1024.8079, 1024.739, 1024.6803, 1024.6575, 1024.5719, 1024.521, NaN, NaN, 1028.6047, 1028.594, 1028.5765, 1028.5533, 1028.5253, 1028.495, 1028.4615, 1028.4148, 1028.3915, 1028.3652, 1028.3298, 1028.2911, 1028.2574, 1028.2274, 1028.1923, 1028.1581, 1028.1095, 1028.0753, 1028.0482, 1028.0159, 1027.9775, 1027.941, 1027.9084, 1027.8683, 1027.832, 1027.7968, 1027.7646, 1027.7361, 1027.7054, 1027.6744, 1027.6392, 1027.6023, 1027.5618, 1027.5286, 1027.4927, 1027.4484, 1027.4, 1027.3551, 1027.3081, 1027.2803, 1027.2501, 1027.2166, 1027.1823, 1027.1484, 1027.1031, 1027.059, 1027.0244, 1026.9873, 1026.9371, 1026.8932, 1026.8539, 1026.8135, 1026.7501, 1026.6973, 1026.6239, 1026.5469, 1026.4734, 1026.386, 1026.3047, 1026.2264, 1026.1602, 1026.0977, 1026.0432, 1025.9763, 1025.8992, 1025.8118, 1025.733, 1025.6194, 1025.501, 1025.3427, 1025.2703, 1025.1942, 1025.067, 1024.8926, 1024.7853, 1024.7407, 1024.675, 1024.5748, 1024.5265, 1024.4546, 1024.4364, NaN, NaN, 1028.5603, 1028.546, 1028.5306, 1028.5123, 1028.4801, 1028.4509, 1028.4182, 1028.3804, 1028.3433, 1028.295, 1028.2609, 1028.233, 1028.2072, 1028.1829, 1028.1569, 1028.128, 1028.0958, 1028.0682, 1028.0336, 1028.0038, 1027.9614, 1027.9269, 1027.89, 1027.8582, 1027.8252, 1027.7927, 1027.7677, 1027.7426, 1027.7141, 1027.6871, 1027.6593, 1027.6276, 1027.6039, 1027.5756, 1027.5402, 1027.5133, 1027.4841, 1027.4454, 1027.4132, 1027.3718, 1027.3336, 1027.3004, 1027.2714, 1027.2332, 1027.1943, 1027.1592, 1027.1184, 1027.0787, 1027.0289, 1026.9858, 1026.9276, 1026.8779, 1026.8228, 1026.774, 1026.7278, 1026.6735, 1026.6185, 1026.545, 1026.4961, 1026.4159, 1026.3499, 1026.2976, 1026.2611, 1026.1974, 1026.0911, 1025.9772, 1025.8995, 1025.8146, 1025.73, 1025.6555, 1025.5591, 1025.4623, 1025.3829, 1025.3182, 1025.2107, 1025.0936, 1025.0338, 1024.9032, 1024.7957, 1024.6741, 1024.5511, 1024.4657, 1024.3904, 1024.3619, NaN, NaN, 1028.5607, 1028.5466, 1028.5288, 1028.5106, 1028.484, 1028.4553, 1028.4282, 1028.3925, 1028.361, 1028.3324, 1028.2987, 1028.2584, 1028.2305, 1028.2017, 1028.1655, 1028.1213, 1028.0859, 1028.0549, 1028.0193, 1027.9729, 1027.9381, 1027.9005, 1027.8651, 1027.833, 1027.8024, 1027.7706, 1027.7374, 1027.7052, 1027.673, 1027.6394, 1027.6046, 1027.5752, 1027.5408, 1027.5044, 1027.4741, 1027.4325, 1027.3911, 1027.3391, 1027.2943, 1027.2614, 1027.2312, 1027.2006, 1027.1627, 1027.1285, 1027.1017, 1027.0648, 1027.0267, 1026.9769, 1026.9286, 1026.8605, 1026.8116, 1026.7653, 1026.6987, 1026.62, 1026.5281, 1026.4149, 1026.3549, 1026.3079, 1026.2695, 1026.1666, 1026.0615, 1025.9576, 1025.8748, 1025.752, 1025.6573, 1025.5437, 1025.4581, 1025.3701, 1025.2758, 1025.2112, 1025.1409, 1025.055, 1024.9619, 1024.8906, 1024.8524, 1024.7695, 1024.6819, 1024.5753, 1024.4362, 1024.3737, NaN, NaN, 1028.6193, 1028.6064, 1028.5847, 1028.5518, 1028.516, 1028.4858, 1028.4481, 1028.418, 1028.3894, 1028.3508, 1028.3175, 1028.2927, 1028.2684, 1028.2405, 1028.2126, 1028.184, 1028.15, 1028.1233, 1028.095, 1028.0654, 1028.0269, 1027.993, 1027.9622, 1027.9314, 1027.8896, 1027.8566, 1027.8235, 1027.7899, 1027.7606, 1027.7351, 1027.7078, 1027.6838, 1027.657, 1027.625, 1027.5955, 1027.5662, 1027.5304, 1027.5043, 1027.4833, 1027.453, 1027.4142, 1027.3853, 1027.3566, 1027.3237, 1027.2869, 1027.2499, 1027.2151, 1027.1866, 1027.1558, 1027.1288, 1027.1018, 1027.0596, 1027.0231, 1026.995, 1026.9592, 1026.9232, 1026.8788, 1026.8378, 1026.7928, 1026.7328, 1026.6603, 1026.5911, 1026.5175, 1026.4237, 1026.3258, 1026.2373, 1026.1482, 1026.0671, 1026.0101, 1025.9136, 1025.8201, 1025.7069, 1025.5697, 1025.489, 1025.3988, 1025.3151, 1025.1565, 1025.0596, 1025.0133, 1024.9607, 1024.9137, 1024.8379, 1024.7472, 1024.6188, 1024.4849, 1024.4078, 1024.3824, 1024.3654, 1024.3562, NaN, NaN, 1028.5919, 1028.5725, 1028.5487, 1028.5165, 1028.4874, 1028.461, 1028.433, 1028.4038, 1028.3678, 1028.3346, 1028.3008, 1028.2601, 1028.2235, 1028.1903, 1028.1484, 1028.1091, 1028.0824, 1028.0573, 1028.0308, 1027.9883, 1027.9492, 1027.9182, 1027.8783, 1027.8413, 1027.8105, 1027.7714, 1027.7444, 1027.71, 1027.6729, 1027.6332, 1027.5945, 1027.5485, 1027.526, 1027.5042, 1027.4731, 1027.4447, 1027.4049, 1027.3682, 1027.3416, 1027.3141, 1027.2899, 1027.2632, 1027.2382, 1027.2146, 1027.192, 1027.1615, 1027.1279, 1027.1072, 1027.0702, 1027.0334, 1026.9913, 1026.9495, 1026.9177, 1026.88, 1026.8207, 1026.7681, 1026.72, 1026.6836, 1026.635, 1026.5728, 1026.5026, 1026.4473, 1026.3654, 1026.3057, 1026.2408, 1026.1719, 1026.1328, 1026.0809, 1026.0374, 1025.9906, 1025.9459, 1025.9142, 1025.8556, 1025.7842, 1025.6938, 1025.5596, 1025.4698, 1025.3678, 1025.2688, 1025.1434, 1025.0046, 1024.9573, 1024.8812, 1024.791, 1024.6538, 1024.5, 1024.331, 1024.3077, NaN, NaN, 1028.477, 1028.46, 1028.4198, 1028.382, 1028.35, 1028.314, 1028.2643, 1028.1749, 1028.1305, 1028.1035, 1028.0768, 1028.0511, 1028.0247, 1027.9973, 1027.9615, 1027.9269, 1027.8944, 1027.8622, 1027.8264, 1027.7872, 1027.7473, 1027.7012, 1027.6602, 1027.6294, 1027.5916, 1027.54, 1027.4922, 1027.4385, 1027.4092, 1027.3691, 1027.3326, 1027.3016, 1027.2804, 1027.2565, 1027.2258, 1027.1837, 1027.1422, 1027.1038, 1027.0701, 1027.0377, 1027.0037, 1026.954, 1026.9065, 1026.8757, 1026.8143, 1026.7518, 1026.6886, 1026.6448, 1026.5575, 1026.4974, 1026.4504, 1026.3835, 1026.294, 1026.1718, 1026.0828, 1026.0531, 1025.9923, 1025.8838, 1025.8307, 1025.7412, 1025.6455, 1025.4794, 1025.3771, 1025.2194, 1025.1161, 1025.0157, 1024.9089, 1024.7885, 1024.638, 1024.4421, 1024.2537, NaN, NaN, 1027.9646, 1027.9398, 1027.9078, 1027.8359, 1027.7776, 1027.7128, 1027.6567, 1027.5953, 1027.5282, 1027.4631, 1027.3975, 1027.3507, 1027.3014, 1027.2468, 1027.1907, 1027.1417, 1027.0989, 1027.057, 1027.0148, 1026.9742, 1026.9249, 1026.8678, 1026.7875, 1026.7383, 1026.6952, 1026.5906, 1026.4701, 1026.3904, 1026.3485, 1026.2717, 1026.195, 1026.0723, 1026.0094, 1025.9128, 1025.7736, 1025.6157, 1025.4641, 1025.306, 1025.1388, 1025.0232, 1024.9147, 1024.8306, 1024.7119, 1024.514, NaN, NaN, 1027.499, 1027.4576, 1027.4081, 1027.3478, 1027.2965, 1027.2478, 1027.2051, 1027.1575, 1027.1102, 1027.0605, 1027.0116, 1026.9705, 1026.9305, 1026.8613, 1026.7694, 1026.7196, 1026.6709, 1026.573, 1026.4149, 1026.2778, 1026.1533, 1025.9233, 1025.7184, 1025.5076, 1025.3672, 1025.2623, 1025.1251, 1024.9685, 1024.8995, 1024.7935, 1024.5994, NaN, NaN, 1027.2521, 1027.2175, 1027.181, 1027.1348, 1027.0908, 1027.0488, 1027.0027, 1026.952, 1026.9045, 1026.8517, 1026.7699, 1026.6844, 1026.5919, 1026.4868, 1026.3865, 1026.2417, 1026.1233, 1025.9672, 1025.749, 1025.5598, 1025.3942, 1025.2606, 1025.1183, 1024.9567, 1024.8749, 1024.8246, 1024.6593, 1024.4606, NaN, NaN, 1027.1559, 1027.1345, 1027.1073, 1027.0637, 1027.0187, 1026.9607, 1026.9131, 1026.8629, 1026.8116, 1026.7196, 1026.631, 1026.5516, 1026.4396, 1026.3208, 1026.1656, 1026.0405, 1025.7784, 1025.5769, 1025.4006, 1025.1927, 1025.0829, 1024.9789, 1024.8848, 1024.7855, 1024.6093, NaN, NaN, 1027.1421, 1027.1226, 1027.096, 1027.0568, 1027.007, 1026.9586, 1026.9061, 1026.8545, 1026.8005, 1026.7306, 1026.6487, 1026.5625, 1026.4344, 1026.2963, 1026.1078, 1025.8645, 1025.5289, 1025.3296, 1025.166, 1025.0596, 1024.8953, 1024.7832, 1024.6124, NaN, NaN, 1027.1277, 1027.1063, 1027.0751, 1027.0325, 1026.9875, 1026.9359, 1026.8779, 1026.8131, 1026.7373, 1026.6528, 1026.5778, 1026.5328, 1026.4553, 1026.3756, 1026.237, 1026.0365, 1025.7734, 1025.5941, 1025.4655, 1025.3025, 1025.1987, 1025.09, 1024.8892, 1024.732, 1024.6407, NaN, NaN, 1027.0775, 1027.0564, 1027.0283, 1026.9882, 1026.942, 1026.8975, 1026.834, 1026.765, 1026.6805, 1026.5912, 1026.4283, 1026.2783, 1026.1276, 1025.9568, 1025.6718, 1025.4717, 1025.3021, 1025.2561, 1025.216, 1025.0908, 1024.8722, 1024.6597, NaN, NaN, 1027.0593, 1027.038, 1027.0089, 1026.9644, 1026.9176, 1026.8666, 1026.8181, 1026.7566, 1026.6498, 1026.5502, 1026.4081, 1026.2678, 1026.1211, 1025.9221, 1025.6573, 1025.477, 1025.38, 1025.3401, 1025.3035, 1025.1697, 1025.0759, 1024.9292, 1024.7377, 1024.4865, NaN, NaN, 1027.0248, 1027.0052, 1026.978, 1026.9397, 1026.9012, 1026.8593, 1026.8146, 1026.7725, 1026.7175, 1026.6124, 1026.5162, 1026.3903, 1026.2688, 1026.1478, 1026.0193, 1025.8071, 1025.5927, 1025.5056, 1025.3824, 1025.2762, 1025.1626, 1025.064, 1024.9482, 1024.7955, 1024.5737, NaN, NaN, 1026.9835, 1026.9609, 1026.9353, 1026.8947, 1026.8539, 1026.8027, 1026.736, 1026.6497, 1026.5737, 1026.4636, 1026.3333, 1026.2152, 1026.1309, 1025.9203, 1025.7404, 1025.6128, 1025.535, 1025.4377, 1025.2913, 1025.1646, 1025.0719, 1025.0111, 1024.8577, 1024.587, NaN, NaN, 1026.9392, 1026.9165, 1026.89, 1026.8518, 1026.8059, 1026.7473, 1026.6946, 1026.6086, 1026.508, 1026.4131, 1026.2928, 1026.2164, 1026.1152, 1025.9039, 1025.6959, 1025.5547, 1025.4374, 1025.2714, 1025.1442, 1025.0629, 1024.9005, 1024.7412, 1024.5032, NaN, NaN, 1026.8936, 1026.8704, 1026.8364, 1026.7902, 1026.7369, 1026.6649, 1026.6014, 1026.4866, 1026.3501, 1026.2158, 1026.0897, 1025.8589, 1025.6278, 1025.3304, 1025.0198, 1024.7047, 1024.5457, 1024.4989, 1024.4731, NaN, NaN, 1026.85, 1026.819, 1026.7832, 1026.7334, 1026.6744, 1026.5789, 1026.4421, 1026.3107, 1026.2539, 1026.1617, 1026.12, 1026.0778, 1025.957, 1025.8469, 1025.6545, 1025.5469, 1025.3293, 1025.0576, 1024.7928, 1024.5676, 1024.459, 1024.371, NaN, NaN, 1026.7744, 1026.743, 1026.7095, 1026.6631, 1026.5623, 1026.4458, 1026.3065, 1026.1993, 1026.0944, 1025.9932, 1025.8108, 1025.6024, 1025.329, 1025.0477, 1024.7643, 1024.4626, NaN, NaN, 1026.7423, 1026.7202, 1026.689, 1026.6517, 1026.6077, 1026.5515, 1026.4668, 1026.3116, 1026.2098, 1026.1304, 1025.9956, 1025.8899, 1025.6991, 1025.5332, 1025.1888, 1024.9302, 1024.6046, NaN, NaN, 1026.7031, 1026.6799, 1026.6521, 1026.6072, 1026.5509, 1026.4222, 1026.3271, 1026.2511, 1026.1943, 1026.145, 1026.0237, 1025.9087, 1025.7828, 1025.5917, 1025.3951, 1025.119, 1024.7745, NaN, NaN, 1026.705, 1026.6871, 1026.6582, 1026.6173, 1026.5747, 1026.4841, 1026.3804, 1026.2924, 1026.2124, 1026.1652, 1026.0791, 1025.9929, 1025.8782, 1025.7623, 1025.6129, 1025.4103, 1025.1647, 1024.6862, NaN, NaN, 1026.686, 1026.6675, 1026.6404, 1026.598, 1026.5582, 1026.4543, 1026.3364, 1026.251, 1026.1918, 1026.1187, 1026.0195, 1025.9177, 1025.8252, 1025.7723, 1025.6534, 1025.5377, 1025.449, 1025.2421, 1025.0878, 1024.8066, 1024.5697, NaN, NaN, 1026.6481, 1026.6263, 1026.596, 1026.5541, 1026.5084, 1026.4524, 1026.303, 1026.1895, 1026.0585, 1025.8326, 1025.6432, 1025.4336, 1025.2095, 1024.9679, 1024.5159, NaN, NaN, 1026.6389, 1026.6167, 1026.5863, 1026.5455, 1026.4977, 1026.3347, 1026.2415, 1026.0729, 1025.8822, 1025.7294, 1025.5486, 1025.3889, 1025.2246, 1025.1505, 1024.7932, NaN, NaN, 1026.6265, 1026.6036, 1026.5713, 1026.53, 1026.4653, 1026.3099, 1026.2416, 1026.1151, 1026.0286, 1025.9287, 1025.7279, 1025.4966, 1025.3572, 1025.2212, 1024.9843, NaN, NaN, 1026.6016, 1026.5814, 1026.5508, 1026.5176, 1026.4812, 1026.4414, 1026.3153, 1026.2198, 1026.1403, 1025.9475, 1025.7035, 1025.4833, 1025.3778, 1025.2155, 1025.0757, NaN, NaN, 1026.6067, 1026.5847, 1026.5566, 1026.5181, 1026.4745, 1026.3938, 1026.2635, 1026.2009, 1026.1249, 1025.9683, 1025.8359, 1025.6023, 1025.4718, 1025.3892, 1025.2405, 1025.1589, NaN, NaN, 1026.6078, 1026.5851, 1026.5576, 1026.5195, 1026.4692, 1026.3639, 1026.2937, 1026.2352, 1026.1742, 1025.988, 1025.8711, 1025.745, 1025.558, 1025.4541, 1025.3297, 1025.2124, 1025.1301, NaN, NaN, 1026.6023, 1026.5803, 1026.5529, 1026.5133, 1026.4626, 1026.3562, 1026.2886, 1026.2261, 1026.147, 1025.9816, 1025.8667, 1025.7413, 1025.4758, 1025.3102, 1025.1476, NaN, NaN, 1026.5776, 1026.5552, 1026.522, 1026.4707, 1026.4042, 1026.3422, 1026.2875, 1026.2251, 1026.1685, 1026.026, 1025.8713, 1025.7555, 1025.5182, 1025.3348, 1025.1794, 1025.0626, NaN, NaN, 1026.5673, 1026.5459, 1026.5157, 1026.463, 1026.3711, 1026.2997, 1026.217, 1026.0618, 1025.9073, 1025.7214, 1025.4948, 1025.3524, 1025.2554, 1025.0353, NaN, NaN, 1026.5231, 1026.4976, 1026.4617, 1026.3983, 1026.3344, 1026.2666, 1026.1807, 1026.0646, 1025.9127, 1025.7651, 1025.571, 1025.3566, 1025.093, 1025.0012, NaN, NaN, 1026.5061, 1026.4781, 1026.4482, 1026.4092, 1026.3524, 1026.2972, 1026.2069, 1026.1384, 1026.0198, 1025.9083, 1025.8064, 1025.6227, 1025.4441, 1025.2792, 1025.131, 1025.004, NaN, NaN, 1026.4906, 1026.4678, 1026.4365, 1026.3839, 1026.3282, 1026.2645, 1026.1687, 1025.9779, 1025.8184, 1025.618, 1025.4167, 1025.266, 1025.0934, 1025.0302, NaN, NaN, 1026.463, 1026.4413, 1026.4102, 1026.3651, 1026.3108, 1026.2473, 1026.172, 1026.0015, 1025.8551, 1025.7234, 1025.4188, 1025.2375, 1025.1118, 1025.0272, NaN, NaN, 1026.4364, 1026.4143, 1026.3801, 1026.3378, 1026.2936, 1026.2161, 1026.1267, 1026.0276, 1025.8627, 1025.728, 1025.5996, 1025.3018, 1025.1528, 1025.0214, NaN, NaN, 1026.4474, 1026.4193, 1026.3893, 1026.3469, 1026.3142, 1026.2479, 1026.183, 1026.1039, 1025.9548, 1025.8365, 1025.6764, 1025.4872, 1025.2312, 1025.0553, 1025.0062, NaN, NaN, 1026.4094, 1026.3842, 1026.3523, 1026.3135, 1026.269, 1026.2001, 1026.1149, 1026.022, 1025.9164, 1025.8118, 1025.6157, 1025.3074, 1025.0662, 1025.0022, NaN, NaN, 1026.3817, 1026.3604, 1026.3346, 1026.2999, 1026.2572, 1026.185, 1026.115, 1026.0443, 1025.9354, 1025.8485, 1025.7207, 1025.5298, 1025.3375, 1025.1288, 1025.0098, NaN, NaN, 1026.3766, 1026.355, 1026.3221, 1026.2775, 1026.2268, 1026.171, 1026.1239, 1026.0309, 1025.9055, 1025.7286, 1025.5612, 1025.304, 1025.0603, 1024.9935, NaN, NaN, 1026.349, 1026.3251, 1026.2828, 1026.2164, 1026.1656, 1026.1035, 1025.9965, 1025.8588, 1025.6714, 1025.49, 1025.2744, 1025.1227, 1025.0386, 1024.9962, NaN, NaN, 1026.3647, 1026.3298, 1026.267, 1026.2158, 1026.1664, 1026.1047, 1026.0277, 1025.9131, 1025.7623, 1025.625, 1025.5566, 1025.3438, 1025.1855, 1025.0336, NaN, NaN, 1026.2997, 1026.268, 1026.2307, 1026.1843, 1026.1396, 1026.0734, 1026.0114, 1025.9329, 1025.8142, 1025.5743, 1025.3623, 1025.1318, 1025.0372, 1025.017, 1025.0131, NaN, NaN, 1026.2904, 1026.2563, 1026.209, 1026.1564, 1026.112, 1026.0476, 1025.9396, 1025.8344, 1025.6355, 1025.358, 1025.0812, 1024.9647, NaN, NaN, 1026.2532, 1026.2258, 1026.1975, 1026.1544, 1026.1179, 1026.0614, 1025.9789, 1025.8723, 1025.6921, 1025.4048, 1025.221, 1025.0674, 1025.0358, 1025.0243, NaN, NaN, 1026.2806, 1026.2343, 1026.1975, 1026.1537, 1026.0989, 1026.0374, 1025.9441, 1025.8158, 1025.637, 1025.3606, 1025.0781, 1024.9879, NaN, NaN, 1026.2701, 1026.2391, 1026.204, 1026.171, 1026.1311, 1026.0917, 1026.046, 1025.9884, 1025.9142, 1025.8202, 1025.7064, 1025.5205, 1025.3109, 1025.144, 1025.0807, NaN, NaN, 1026.221, 1026.1931, 1026.1544, 1026.1014, 1026.0516, 1025.9877, 1025.8766, 1025.7397, 1025.5602, 1025.2361, 1025.0026, NaN, NaN, 1026.2388, 1026.2139, 1026.1779, 1026.1317, 1026.0858, 1026.0359, 1025.9757, 1025.8823, 1025.7593, 1025.5387, 1025.2102, 1025.0406, 1025.0126, 1025.0135, NaN, NaN, 1026.2095, 1026.1869, 1026.1554, 1026.1086, 1026.0564, 1026.0066, 1025.9297, 1025.7834, 1025.5688, 1025.1978, 1024.9768, NaN, NaN, 1026.2157, 1026.1927, 1026.1594, 1026.1189, 1026.0732, 1026.0093, 1025.9153, 1025.786, 1025.6064, 1025.297, 1025.0924, 1024.9996, 1024.9526, NaN, NaN, 1026.2561, 1026.228, 1026.195, 1026.155, 1026.1139, 1026.058, 1025.987, 1025.873, 1025.7365, 1025.4968, 1025.3059, 1025.1075, 1024.9744, NaN, NaN, 1026.2943, 1026.271, 1026.2369, 1026.1881, 1026.1498, 1026.1007, 1026.0156, 1025.8461, 1025.6813, 1025.4933, 1025.308, 1025.1145, 1024.9993, 1024.9543, NaN, NaN, 1026.2988, 1026.2747, 1026.2473, 1026.2094, 1026.1671, 1026.1178, 1026.0631, 1025.9203, 1025.7451, 1025.504, 1025.2428, 1025.0485, 1024.9872, NaN, NaN, 1026.3517, 1026.3252, 1026.2845, 1026.2391, 1026.1953, 1026.1377, 1026.0621, 1025.9646, 1025.8203, 1025.5543, 1025.2515, 1025.1536, 1025.0564, 1024.9855, 1024.9766, NaN, NaN, 1026.3351, 1026.3003, 1026.2673, 1026.215, 1026.1205, 1026.002, 1025.8888, 1025.7806, 1025.6694, 1025.5698, 1025.295, 1024.996, NaN, NaN, 1026.3921, 1026.3687, 1026.3298, 1026.2865, 1026.2445, 1026.2047, 1026.1439, 1026.0214, 1025.8729, 1025.7566, 1025.6566, 1025.4373, 1025.0936, 1024.9763, NaN, NaN, 1026.4154, 1026.3918, 1026.366, 1026.3258, 1026.287, 1026.2482, 1026.1848, 1026.1248, 1026.0046, 1025.8677, 1025.7491, 1025.634, 1025.396, 1025.1229, 1024.9811, NaN, NaN, 1026.4193, 1026.3978, 1026.3713, 1026.3326, 1026.2872, 1026.2198, 1026.1202, 1025.9722, 1025.8368, 1025.7157, 1025.5581, 1025.389, 1025.2139, 1025.0664, 1024.9504, NaN, NaN, 1026.4296, 1026.3972, 1026.3654, 1026.326, 1026.2891, 1026.2468, 1026.1401, 1026.0372, 1025.9089, 1025.7731, 1025.5623, 1025.3131, 1025.0889, 1024.9324, NaN, NaN, 1026.4907, 1026.4492, 1026.4113, 1026.3663, 1026.3286, 1026.2924, 1026.1962, 1026.1028, 1026.0076, 1025.8972, 1025.7737, 1025.6542, 1025.4346, 1025.1044, NaN, NaN, 1026.5527, 1026.5253, 1026.4778, 1026.4264, 1026.3627, 1026.3054, 1026.2152, 1026.1143, 1025.9905, 1025.8896, 1025.7599, 1025.6489, 1025.4949, 1025.2095, 1024.9714, NaN, NaN, 1026.5856, 1026.5614, 1026.5261, 1026.4741, 1026.3773, 1026.2825, 1026.2059, 1026.1426, 1026.0385, 1025.9204, 1025.7847, 1025.6395, 1025.4388, 1025.1526, 1024.9785, NaN, NaN, 1026.6313, 1026.6107, 1026.5854, 1026.551, 1026.4728, 1026.3726, 1026.2943, 1026.2222, 1026.1067, 1025.9645, 1025.8356, 1025.6724, 1025.4818, 1025.3868, 1025.2836, 1025.1412, 1025.003, NaN, NaN, 1026.6185, 1026.5974, 1026.5712, 1026.5332, 1026.4481, 1026.3741, 1026.2933, 1026.1943, 1026.106, 1025.9885, 1025.8572, 1025.7278, 1025.559, 1025.4166, 1025.2175, 1025.1256, 1024.9863, NaN, NaN, 1026.6613, 1026.6375, 1026.6074, 1026.5237, 1026.4393, 1026.3661, 1026.2831, 1026.1859, 1026.0491, 1025.922, 1025.7562, 1025.6329, 1025.4166, 1025.1642, 1025.0293, 1024.9601, NaN, NaN, 1026.6781, 1026.6573, 1026.6255, 1026.552, 1026.4565, 1026.3951, 1026.3151, 1026.2485, 1026.146, 1026.0004, 1025.8978, 1025.7543, 1025.5768, 1025.3608, 1025.1989, 1024.9254, NaN, NaN, 1026.6836, 1026.6571, 1026.6056, 1026.5106, 1026.4371, 1026.3374, 1026.2554, 1026.1625, 1026.0203, 1025.8882, 1025.7491, 1025.5957, 1025.4272, 1025.2808, 1025.0536, 1024.8853, NaN, NaN, 1026.6954, 1026.6744, 1026.6469, 1026.5758, 1026.4844, 1026.3864, 1026.3007, 1026.2184, 1026.1342, 1026.0322, 1025.8763, 1025.7468, 1025.5863, 1025.479, 1025.3192, 1025.1917, 1024.9531, NaN, NaN, 1026.7117, 1026.69, 1026.6587, 1026.5978, 1026.4956, 1026.3976, 1026.2902, 1026.2263, 1026.1486, 1026.0494, 1025.8744, 1025.7008, 1025.4604, 1025.2877, 1025.2085, 1025.0648, 1024.9227, NaN, NaN, 1026.7203, 1026.6908, 1026.6414, 1026.5677, 1026.4658, 1026.3687, 1026.2993, 1026.2405, 1026.1605, 1026.0768, 1026.004, 1025.9088, 1025.7386, 1025.4896, 1025.2869, 1025.1442, 1024.9015, NaN, NaN, 1026.7539, 1026.7333, 1026.706, 1026.6216, 1026.5292, 1026.4459, 1026.3881, 1026.3127, 1026.2406, 1026.1746, 1026.1143, 1026.0428, 1025.9158, 1025.7025, 1025.4525, 1025.2723, 1025.1667, 1024.952, 1024.796, NaN, NaN, 1026.7692, 1026.7443, 1026.6935, 1026.6389, 1026.5851, 1026.5146, 1026.426, 1026.359, 1026.2733, 1026.1998, 1026.0862, 1025.9778, 1025.7987, 1025.6157, 1025.4366, 1025.2877, 1025.1962, 1024.8964, 1024.7783, NaN, NaN, 1026.7878, 1026.7635, 1026.6815, 1026.5876, 1026.5135, 1026.4188, 1026.3268, 1026.2445, 1026.1454, 1026.0088, 1025.8981, 1025.7875, 1025.6302, 1025.4021, 1025.2783, 1025.0607, 1024.816, 1024.7247, NaN, NaN, 1026.8073, 1026.7885, 1026.7598, 1026.6932, 1026.5992, 1026.5387, 1026.4669, 1026.3961, 1026.3011, 1026.2019, 1026.0737, 1025.9127, 1025.7804, 1025.5907, 1025.417, 1025.3027, 1025.1547, 1025.046, 1024.7141, 1024.569, NaN, NaN, 1026.8939, 1026.8706, 1026.8379, 1026.8003, 1026.7437, 1026.6351, 1026.5588, 1026.4996, 1026.452, 1026.3566, 1026.2545, 1026.1802, 1026.0537, 1025.9387, 1025.7736, 1025.6482, 1025.5033, 1025.3707, 1025.2593, 1025.1263, 1024.8922, 1024.6272, 1024.5231, NaN, NaN, 1026.9546, 1026.9233, 1026.8875, 1026.8208, 1026.7494, 1026.6594, 1026.5884, 1026.5272, 1026.4564, 1026.3931, 1026.2899, 1026.1774, 1026.0272, 1025.9167, 1025.8009, 1025.612, 1025.407, 1025.2769, 1025.1089, 1024.945, 1024.5677, 1024.4609, NaN, NaN, 1027.0132, 1026.9753, 1026.9171, 1026.8413, 1026.7814, 1026.705, 1026.6384, 1026.5535, 1026.4755, 1026.4071, 1026.3433, 1026.2487, 1026.1774, 1026.0731, 1025.9209, 1025.8018, 1025.5892, 1025.3776, 1025.2152, 1025.1077, 1024.9049, 1024.6892, 1024.4851, NaN, NaN, 1027.0613, 1027.0177, 1026.9568, 1026.8876, 1026.831, 1026.765, 1026.6986, 1026.6334, 1026.584, 1026.5095, 1026.4385, 1026.372, 1026.275, 1026.2223, 1026.1212, 1025.9509, 1025.7246, 1025.4257, 1025.25, 1025.0768, 1024.8866, 1024.7395, 1024.464, 1024.3826, NaN, NaN, 1027.0908, 1027.0491, 1026.9878, 1026.8927, 1026.8397, 1026.7761, 1026.7258, 1026.6564, 1026.5828, 1026.5326, 1026.4663, 1026.3984, 1026.3015, 1026.218, 1026.1207, 1025.9918, 1025.848, 1025.6094, 1025.3712, 1025.2113, 1025.0387, 1024.7123, 1024.4052, 1024.3085, 1024.277, NaN, NaN, 1027.1586, 1027.1226, 1027.0632, 1026.9807, 1026.915, 1026.8594, 1026.7736, 1026.7115, 1026.6543, 1026.5642, 1026.4694, 1026.383, 1026.2878, 1026.2058, 1026.0834, 1025.9087, 1025.761, 1025.5906, 1025.3872, 1025.2123, 1025.0541, 1024.6938, 1024.367, 1024.3347, NaN, NaN, 1027.2183, 1027.1824, 1027.139, 1027.0948, 1027.0223, 1026.9629, 1026.8754, 1026.7704, 1026.6897, 1026.6394, 1026.5856, 1026.4977, 1026.4099, 1026.3054, 1026.1967, 1026.089, 1025.9622, 1025.785, 1025.5311, 1025.3292, 1025.2102, 1025.0125, 1024.7026, 1024.4368, 1024.3805, 1024.3636, NaN, NaN, 1027.3121, 1027.284, 1027.2526, 1027.2134, 1027.1718, 1027.0986, 1027.0222, 1026.9387, 1026.8573, 1026.7787, 1026.7142, 1026.6412, 1026.5525, 1026.4529, 1026.3639, 1026.2701, 1026.1571, 1026.0452, 1025.922, 1025.7645, 1025.556, 1025.3896, 1025.2445, 1025.1057, 1024.8274, 1024.475, 1024.3903, 1024.3483, 1024.3315, NaN, NaN, 1027.4805, 1027.4542, 1027.4154, 1027.3528, 1027.2925, 1027.2485, 1027.2029, 1027.1378, 1027.0605, 1026.9596, 1026.895, 1026.8351, 1026.7822, 1026.7297, 1026.6495, 1026.5828, 1026.4801, 1026.4191, 1026.3488, 1026.2532, 1026.1542, 1026.0404, 1025.8593, 1025.6375, 1025.451, 1025.3127, 1025.1807, 1025.0137, 1024.8112, 1024.4521, 1024.3016, 1024.2753, NaN, NaN, 1027.9751, 1027.926, 1027.8672, 1027.8192, 1027.7839, 1027.7471, 1027.7086, 1027.668, 1027.619, 1027.5597, 1027.5037, 1027.4408, 1027.3915, 1027.3418, 1027.274, 1027.2046, 1027.1196, 1027.0364, 1026.9838, 1026.9382, 1026.8591, 1026.7842, 1026.7097, 1026.6245, 1026.5192, 1026.3961, 1026.3167, 1026.2572, 1026.1519, 1025.9624, 1025.7616, 1025.6102, 1025.4635, 1025.3066, 1025.1659, 1024.9961, 1024.8102, 1024.5695, 1024.3246, 1024.2609, 1024.2397, NaN, NaN, 1028.5172, 1028.4813, 1028.4233, 1028.362, 1028.3026, 1028.2361, 1028.1733, 1028.1128, 1028.0645, 1028.0079, 1027.9552, 1027.9052, 1027.858, 1027.8076, 1027.7623, 1027.7094, 1027.6578, 1027.605, 1027.5529, 1027.506, 1027.4573, 1027.3932, 1027.3282, 1027.2782, 1027.2018, 1027.144, 1027.0878, 1027.0253, 1026.9572, 1026.8947, 1026.8328, 1026.7428, 1026.6752, 1026.6135, 1026.5442, 1026.4503, 1026.3633, 1026.2992, 1026.2173, 1026.109, 1025.8889, 1025.7493, 1025.6272, 1025.4415, 1025.2532, 1025.0853, 1024.9023, 1024.6943, 1024.4514, 1024.2455, 1024.2083, 1024.183, NaN, NaN, 1029.1974, 1029.1732, 1029.1444, 1029.0925, 1029.0526, 1028.9994, 1028.9146, 1028.8685, 1028.8324, 1028.7938, 1028.7413, 1028.6945, 1028.6462, 1028.605, 1028.555, 1028.5029, 1028.4473, 1028.4028, 1028.3579, 1028.312, 1028.2526, 1028.2015, 1028.1622, 1028.1185, 1028.0636, 1028.0203, 1027.9818, 1027.9294, 1027.8793, 1027.833, 1027.777, 1027.7213, 1027.6764, 1027.6322, 1027.5854, 1027.5383, 1027.4902, 1027.4475, 1027.393, 1027.3461, 1027.2909, 1027.2255, 1027.1564, 1027.1001, 1027.0408, 1026.9769, 1026.9185, 1026.8618, 1026.8026, 1026.7319, 1026.6624, 1026.5857, 1026.4799, 1026.3787, 1026.3201, 1026.2601, 1026.1707, 1026.0446, 1025.8833, 1025.7301, 1025.5021, 1025.3201, 1025.1902, 1025.0924, 1024.9637, 1024.9061, 1024.7001, 1024.3318, 1024.268, 1024.1968, 1024.1711, NaN, NaN, 1029.2601, 1029.2372, 1029.2023, 1029.1304, 1029.0686, 1029.018, 1028.9652, 1028.9136, 1028.8627, 1028.8076, 1028.7606, 1028.7035, 1028.6521, 1028.6088, 1028.5542, 1028.5089, 1028.4637, 1028.4073, 1028.3595, 1028.3145, 1028.2615, 1028.2074, 1028.1566, 1028.1108, 1028.0609, 1028.0135, 1027.964, 1027.9104, 1027.8616, 1027.8048, 1027.7551, 1027.6989, 1027.6394, 1027.5896, 1027.5477, 1027.4972, 1027.45, 1027.3922, 1027.3453, 1027.2922, 1027.2322, 1027.1809, 1027.1185, 1027.0543, 1026.9966, 1026.923, 1026.8522, 1026.7894, 1026.714, 1026.657, 1026.5758, 1026.4735, 1026.3746, 1026.2509, 1026.1406, 1025.9481, 1025.7468, 1025.6328, 1025.5208, 1025.3916, 1025.2494, 1025.1199, 1024.9487, 1024.7578, 1024.446, 1024.3164, 1024.2136, 1024.1665, 1024.1311, NaN, NaN, 1029.2351, 1029.2112, 1029.1776, 1029.1311, 1029.091, 1029.0454, 1028.9978, 1028.9485, 1028.9015, 1028.8503, 1028.7988, 1028.7476, 1028.7013, 1028.6539, 1028.6042, 1028.5483, 1028.497, 1028.4515, 1028.4061, 1028.3639, 1028.311, 1028.2584, 1028.2015, 1028.1582, 1028.1141, 1028.0665, 1028.0221, 1027.974, 1027.9283, 1027.8826, 1027.8276, 1027.7826, 1027.7329, 1027.6793, 1027.6278, 1027.5781, 1027.5304, 1027.4794, 1027.4266, 1027.371, 1027.3109, 1027.2633, 1027.1938, 1027.1227, 1027.0524, 1026.9697, 1026.8995, 1026.8252, 1026.742, 1026.6433, 1026.532, 1026.4384, 1026.3206, 1026.2336, 1026.1211, 1026.0026, 1025.8961, 1025.7408, 1025.5912, 1025.5127, 1025.388, 1025.2946, 1025.1508, 1025.0151, 1024.9213, 1024.7733, 1024.5654, 1024.4319, 1024.2787, 1024.1869, 1024.1357, 1024.0874, NaN, NaN, 1029.2283, 1029.2001, 1029.1655, 1029.121, 1029.077, 1029.0306, 1028.9849, 1028.9407, 1028.899, 1028.852, 1028.8124, 1028.7734, 1028.7299, 1028.6863, 1028.6437, 1028.5975, 1028.5499, 1028.5017, 1028.4602, 1028.4224, 1028.3712, 1028.3192, 1028.2712, 1028.2291, 1028.1783, 1028.1257, 1028.0782, 1028.0295, 1027.9818, 1027.934, 1027.8849, 1027.8407, 1027.7922, 1027.7427, 1027.6948, 1027.6459, 1027.5903, 1027.5297, 1027.477, 1027.4213, 1027.368, 1027.3104, 1027.2563, 1027.1868, 1027.1185, 1027.0566, 1027.0056, 1026.919, 1026.8164, 1026.7263, 1026.6614, 1026.5905, 1026.4697, 1026.3295, 1026.192, 1026.0994, 1025.9463, 1025.8127, 1025.6165, 1025.4922, 1025.3754, 1025.2708, 1025.0996, 1024.9071, 1024.7278, 1024.5309, 1024.423, 1024.2972, 1024.186, 1024.1283, 1024.0621, 1024.0056, NaN, NaN, 1029.2344, 1029.1985, 1029.1593, 1029.1144, 1029.0802, 1029.0342, 1028.989, 1028.9482, 1028.9045, 1028.8613, 1028.82, 1028.7714, 1028.7274, 1028.6855, 1028.6422, 1028.5956, 1028.5482, 1028.4957, 1028.4556, 1028.4025, 1028.3579, 1028.3103, 1028.2656, 1028.2217, 1028.1774, 1028.1296, 1028.0824, 1028.0355, 1027.9893, 1027.9426, 1027.8912, 1027.845, 1027.7947, 1027.7448, 1027.6982, 1027.6488, 1027.5946, 1027.5488, 1027.5043, 1027.4532, 1027.4003, 1027.3469, 1027.2999, 1027.249, 1027.1843, 1027.1205, 1027.0525, 1026.9698, 1026.8994, 1026.8256, 1026.7194, 1026.6504, 1026.5283, 1026.4199, 1026.3055, 1026.1542, 1026.0138, 1025.8606, 1025.7196, 1025.5819, 1025.4495, 1025.3407, 1025.2683, 1025.1672, 1024.9886, 1024.7601, 1024.5887, 1024.4402, 1024.3188, 1024.1821, 1024.0852, 1024.0623, NaN, NaN, 1029.222, 1029.1947, 1029.1564, 1029.1122, 1029.0593, 1029.0089, 1028.9688, 1028.9187, 1028.8735, 1028.821, 1028.7703, 1028.7198, 1028.6648, 1028.6154, 1028.5713, 1028.5159, 1028.4629, 1028.4171, 1028.3684, 1028.3214, 1028.2654, 1028.21, 1028.1647, 1028.1158, 1028.0712, 1028.025, 1027.9733, 1027.9227, 1027.8652, 1027.812, 1027.7651, 1027.7157, 1027.6636, 1027.6107, 1027.5562, 1027.5051, 1027.4501, 1027.3987, 1027.3507, 1027.3036, 1027.2512, 1027.1924, 1027.123, 1027.051, 1026.9749, 1026.889, 1026.8176, 1026.7117, 1026.6279, 1026.5002, 1026.369, 1026.238, 1026.0549, 1025.919, 1025.8141, 1025.6993, 1025.569, 1025.4188, 1025.3148, 1025.2197, 1025.1053, 1024.9802, 1024.8154, 1024.6385, 1024.4585, 1024.4089, 1024.3346, 1024.2357, 1024.1493, 1024.0715, 1024.051, NaN, NaN, 1029.2266, 1029.198, 1029.1676, 1029.1218, 1029.0781, 1029.0378, 1028.9973, 1028.9529, 1028.9075, 1028.8613, 1028.8114, 1028.7662, 1028.7191, 1028.6698, 1028.6195, 1028.5735, 1028.5222, 1028.4802, 1028.4337, 1028.3824, 1028.3263, 1028.2755, 1028.2338, 1028.1805, 1028.1285, 1028.0798, 1028.0271, 1027.9705, 1027.9159, 1027.8638, 1027.8159, 1027.7626, 1027.7103, 1027.6512, 1027.5975, 1027.547, 1027.4972, 1027.4462, 1027.3943, 1027.3291, 1027.2699, 1027.1982, 1027.1273, 1027.0569, 1026.9917, 1026.9159, 1026.8394, 1026.7422, 1026.6501, 1026.5377, 1026.419, 1026.2859, 1026.1488, 1025.9697, 1025.8092, 1025.6616, 1025.497, 1025.3849, 1025.2883, 1025.2052, 1025.0636, 1024.8611, 1024.7098, 1024.5427, 1024.3912, 1024.2349, 1024.0924, 1024.0248, 1023.98224, 1023.9554, NaN, NaN, 1029.2301, 1029.203, 1029.1672, 1029.1184, 1029.0709, 1029.0244, 1028.9767, 1028.9358, 1028.8912, 1028.8458, 1028.7977, 1028.7545, 1028.7069, 1028.6598, 1028.6165, 1028.5713, 1028.526, 1028.4758, 1028.4333, 1028.3931, 1028.3502, 1028.2976, 1028.2478, 1028.1979, 1028.1539, 1028.1003, 1028.0486, 1027.9974, 1027.9453, 1027.8945, 1027.8337, 1027.7869, 1027.7434, 1027.6952, 1027.6416, 1027.596, 1027.5431, 1027.4904, 1027.4385, 1027.3878, 1027.3317, 1027.2642, 1027.2092, 1027.1511, 1027.0894, 1027.0116, 1026.9354, 1026.8529, 1026.7931, 1026.7148, 1026.6151, 1026.509, 1026.407, 1026.3065, 1026.1417, 1025.9598, 1025.8394, 1025.7233, 1025.5868, 1025.4388, 1025.294, 1025.147, 1025.0262, 1024.8434, 1024.7173, 1024.5869, 1024.449, 1024.3151, 1024.1415, 1023.93713, 1023.8898, 1023.8521, 1023.822, 1023.8052, NaN, NaN, 1029.2339, 1029.2081, 1029.172, 1029.1296, 1029.0857, 1029.042, 1028.9988, 1028.9532, 1028.9132, 1028.8705, 1028.8271, 1028.781, 1028.7385, 1028.6907, 1028.6467, 1028.6078, 1028.5654, 1028.5254, 1028.4791, 1028.4363, 1028.3949, 1028.3519, 1028.3083, 1028.2673, 1028.2242, 1028.1793, 1028.1356, 1028.0901, 1028.0458, 1028.0052, 1027.9631, 1027.9137, 1027.8711, 1027.8209, 1027.7784, 1027.7345, 1027.6923, 1027.6453, 1027.5975, 1027.5576, 1027.5094, 1027.4653, 1027.4174, 1027.3674, 1027.3131, 1027.2446, 1027.1865, 1027.1311, 1027.064, 1027.0065, 1026.9369, 1026.8579, 1026.7826, 1026.7156, 1026.6167, 1026.4829, 1026.3938, 1026.2421, 1026.119, 1025.976, 1025.7875, 1025.6549, 1025.5297, 1025.3895, 1025.2804, 1025.1769, 1025.0815, 1024.9884, 1024.8019, 1024.5925, 1024.3617, 1024.1888, 1024.1005, 1023.9642, 1023.821, 1023.7919, 1023.76855, 1023.7511, NaN, NaN, 1029.2385, 1029.214, 1029.179, 1029.1324, 1029.0916, 1029.0448, 1029.0055, 1028.9633, 1028.922, 1028.8745, 1028.8268, 1028.7793, 1028.7373, 1028.6895, 1028.6445, 1028.6035, 1028.5618, 1028.5112, 1028.4592, 1028.4128, 1028.3694, 1028.3236, 1028.2708, 1028.2227, 1028.1796, 1028.1305, 1028.0886, 1028.045, 1027.9963, 1027.9512, 1027.9056, 1027.8584, 1027.8104, 1027.7682, 1027.7302, 1027.6891, 1027.6425, 1027.5941, 1027.5396, 1027.4808, 1027.4347, 1027.3802, 1027.3248, 1027.2676, 1027.1979, 1027.1299, 1027.0801, 1027.0139, 1026.9315, 1026.8331, 1026.7172, 1026.5975, 1026.464, 1026.3248, 1026.2216, 1026.0945, 1025.9679, 1025.8424, 1025.7052, 1025.6075, 1025.4945, 1025.3668, 1025.2827, 1025.1426, 1024.9799, 1024.8109, 1024.6616, 1024.5653, 1024.3638, 1024.1719, 1024.0807, 1023.9798, 1023.7718, 1023.74725, 1023.7267, 1023.7135, NaN, NaN, 1029.2214, 1029.1962, 1029.1664, 1029.118, 1029.069, 1029.022, 1028.9747, 1028.9287, 1028.8763, 1028.8259, 1028.7803, 1028.7345, 1028.6857, 1028.6375, 1028.5927, 1028.5503, 1028.5051, 1028.4609, 1028.4164, 1028.3656, 1028.3198, 1028.2728, 1028.2275, 1028.1736, 1028.1252, 1028.0715, 1028.0181, 1027.9618, 1027.9137, 1027.8522, 1027.7983, 1027.7448, 1027.6869, 1027.6351, 1027.5836, 1027.5282, 1027.4645, 1027.408, 1027.3499, 1027.2842, 1027.2063, 1027.1489, 1027.085, 1027.0166, 1026.946, 1026.8586, 1026.7736, 1026.6613, 1026.532, 1026.4105, 1026.323, 1026.1902, 1026.0768, 1025.8903, 1025.7467, 1025.622, 1025.511, 1025.3976, 1025.2689, 1025.1202, 1024.9888, 1024.896, 1024.8057, 1024.6554, 1024.5339, 1024.2911, 1024.1129, 1024.036, 1023.78546, 1023.7232, 1023.695, 1023.6808, NaN, NaN, 1029.2211, 1029.1923, 1029.158, 1029.1056, 1029.0575, 1029.0111, 1028.9608, 1028.9177, 1028.8711, 1028.8204, 1028.7701, 1028.7198, 1028.673, 1028.6261, 1028.5825, 1028.5364, 1028.4932, 1028.4469, 1028.3971, 1028.352, 1028.3069, 1028.257, 1028.2017, 1028.1501, 1028.0992, 1028.0476, 1027.9883, 1027.9396, 1027.883, 1027.835, 1027.7806, 1027.7318, 1027.681, 1027.635, 1027.578, 1027.5189, 1027.4633, 1027.4025, 1027.3445, 1027.2798, 1027.2267, 1027.1631, 1027.0984, 1027.0295, 1026.9402, 1026.8525, 1026.756, 1026.6437, 1026.4587, 1026.3318, 1026.1285, 1025.9928, 1025.8862, 1025.7631, 1025.6504, 1025.5161, 1025.4098, 1025.2721, 1025.1312, 1025.0182, 1024.9425, 1024.808, 1024.6847, 1024.5369, 1024.3848, 1024.2234, 1024.0924, 1024.0421, 1023.9, 1023.65686, 1023.6337, 1023.6178, NaN, NaN, 1029.2391, 1029.2146, 1029.1788, 1029.1292, 1029.0773, 1029.0216, 1028.9634, 1028.9172, 1028.8683, 1028.8182, 1028.771, 1028.7212, 1028.6741, 1028.6238, 1028.5703, 1028.5168, 1028.4667, 1028.4194, 1028.369, 1028.3173, 1028.2694, 1028.2189, 1028.1753, 1028.1261, 1028.0742, 1028.0275, 1027.9777, 1027.9253, 1027.8705, 1027.8231, 1027.7751, 1027.7242, 1027.673, 1027.6252, 1027.5778, 1027.5299, 1027.4791, 1027.4227, 1027.3671, 1027.3093, 1027.2354, 1027.161, 1027.0969, 1027.0237, 1026.9388, 1026.8435, 1026.7648, 1026.6492, 1026.5436, 1026.4607, 1026.358, 1026.1881, 1026.031, 1025.8767, 1025.7513, 1025.5924, 1025.4569, 1025.3464, 1025.236, 1025.0924, 1025.0106, 1024.8789, 1024.7561, 1024.5931, 1024.4032, 1024.263, 1024.1039, 1024.0186, 1023.744, 1023.6531, 1023.62726, 1023.6097, NaN, NaN, 1029.2307, 1029.2068, 1029.1732, 1029.1226, 1029.077, 1029.0325, 1028.9867, 1028.9384, 1028.8911, 1028.8424, 1028.7941, 1028.747, 1028.6967, 1028.6486, 1028.601, 1028.5566, 1028.5099, 1028.4578, 1028.4071, 1028.3574, 1028.3115, 1028.2607, 1028.2119, 1028.1625, 1028.1112, 1028.0626, 1028.0139, 1027.9635, 1027.9109, 1027.8588, 1027.8058, 1027.7529, 1027.6941, 1027.6425, 1027.5874, 1027.537, 1027.48, 1027.4232, 1027.3595, 1027.3003, 1027.2323, 1027.1697, 1027.1145, 1027.0547, 1026.9801, 1026.8972, 1026.7959, 1026.7063, 1026.5774, 1026.4714, 1026.3593, 1026.2103, 1026.0232, 1025.8898, 1025.8008, 1025.7023, 1025.5944, 1025.4535, 1025.331, 1025.1969, 1025.1206, 1025.0255, 1024.8998, 1024.7368, 1024.5569, 1024.413, 1024.3203, 1024.2352, 1024.1326, 1024.0576, 1023.83905, 1023.6724, 1023.6484, 1023.632, NaN, NaN, 1029.2314, 1029.2054, 1029.1713, 1029.1311, 1029.0819, 1029.0356, 1028.9852, 1028.9418, 1028.899, 1028.8452, 1028.8043, 1028.7587, 1028.7078, 1028.6564, 1028.61, 1028.564, 1028.5167, 1028.4655, 1028.416, 1028.3668, 1028.3188, 1028.2693, 1028.2168, 1028.1671, 1028.1193, 1028.0751, 1028.0168, 1027.9663, 1027.9178, 1027.8699, 1027.8118, 1027.7579, 1027.7095, 1027.6583, 1027.6012, 1027.5488, 1027.497, 1027.44, 1027.381, 1027.3207, 1027.269, 1027.2083, 1027.1421, 1027.0608, 1026.9805, 1026.9082, 1026.83, 1026.7445, 1026.6575, 1026.5546, 1026.3972, 1026.2594, 1026.1382, 1025.999, 1025.8154, 1025.7169, 1025.6426, 1025.5264, 1025.3876, 1025.2283, 1025.1117, 1025.0187, 1024.8673, 1024.7314, 1024.5272, 1024.4465, 1024.3075, 1024.2213, 1024.1426, 1024.0186, 1023.7096, 1023.66656, 1023.65027, 1023.64, NaN, NaN, 1029.2421, 1029.2156, 1029.177, 1029.1364, 1029.0894, 1029.0417, 1028.9885, 1028.9469, 1028.9037, 1028.8585, 1028.8091, 1028.7607, 1028.713, 1028.6638, 1028.6139, 1028.5618, 1028.5092, 1028.4567, 1028.4059, 1028.3557, 1028.3059, 1028.2578, 1028.2086, 1028.1578, 1028.1056, 1028.0533, 1028.0049, 1027.9596, 1027.9092, 1027.8591, 1027.816, 1027.7653, 1027.7162, 1027.667, 1027.6154, 1027.5598, 1027.5057, 1027.4464, 1027.3945, 1027.3325, 1027.2637, 1027.1929, 1027.1096, 1027.043, 1026.9792, 1026.8961, 1026.8079, 1026.7515, 1026.6451, 1026.5352, 1026.4103, 1026.3047, 1026.1208, 1025.9492, 1025.7726, 1025.6111, 1025.4817, 1025.3147, 1025.2054, 1025.0881, 1024.943, 1024.6875, 1024.5911, 1024.4961, 1024.404, 1024.2968, 1024.1934, 1024.0864, 1023.8632, 1023.6712, 1023.6515, NaN, NaN, 1029.24, 1029.2134, 1029.1805, 1029.1311, 1029.0758, 1029.0228, 1028.9734, 1028.9181, 1028.8646, 1028.8134, 1028.764, 1028.7109, 1028.6582, 1028.6079, 1028.5603, 1028.5001, 1028.4521, 1028.4253, 1028.3683, 1028.3136, 1028.2655, 1028.2131, 1028.1583, 1028.1083, 1028.0537, 1028.003, 1027.9523, 1027.9095, 1027.8545, 1027.8076, 1027.7576, 1027.7065, 1027.6528, 1027.5999, 1027.5464, 1027.4902, 1027.4414, 1027.381, 1027.328, 1027.2672, 1027.21, 1027.1365, 1027.0621, 1026.9838, 1026.9095, 1026.8038, 1026.7054, 1026.6056, 1026.5304, 1026.4045, 1026.2688, 1026.135, 1025.9635, 1025.8038, 1025.6803, 1025.522, 1025.3933, 1025.274, 1025.1082, 1024.9749, 1024.7539, 1024.6156, 1024.5459, 1024.4706, 1024.3507, 1024.2244, 1024.15, 1023.98334, 1023.69275, 1023.6735, 1023.6551, NaN, NaN, 1029.211, 1029.1831, 1029.143, 1029.0955, 1029.0507, 1029.0072, 1028.9641, 1028.9165, 1028.8635, 1028.8104, 1028.7596, 1028.7075, 1028.6603, 1028.6152, 1028.57, 1028.5262, 1028.4753, 1028.4281, 1028.378, 1028.3242, 1028.274, 1028.2224, 1028.1731, 1028.1176, 1028.0635, 1028.0094, 1027.9537, 1027.904, 1027.8477, 1027.7916, 1027.7334, 1027.6768, 1027.6235, 1027.5668, 1027.5164, 1027.4672, 1027.4086, 1027.3436, 1027.2816, 1027.2305, 1027.1707, 1027.0844, 1027.0381, 1027.0205, 1026.95, 1026.5145, 1026.1826, 1026.0109, 1025.9812, 1025.728, 1025.7776, 1026.1726, 1025.8766, 1025.591, 1025.4775, 1025.4221, 1025.282, 1025.1724, 1025.0328, 1024.8673, 1024.7472, 1024.5596, 1024.5063, 1024.447, 1024.3209, 1024.2057, 1024.143, 1023.99866, 1023.70233, 1023.6786, 1023.6674, NaN, NaN, 1029.1951, 1029.168, 1029.1335, 1029.0823, 1029.0308, 1028.972, 1028.9209, 1028.8713, 1028.8174, 1028.765, 1028.7179, 1028.6707, 1028.6211, 1028.5668, 1028.5145, 1028.4629, 1028.4126, 1028.3635, 1028.3176, 1028.269, 1028.2196, 1028.1687, 1028.1172, 1028.0663, 1028.0114, 1027.9591, 1027.9005, 1027.8451, 1027.7925, 1027.7377, 1027.6913, 1027.6351, 1027.5837, 1027.5376, 1027.4885, 1027.4285, 1027.3735, 1027.3168, 1027.2627, 1027.2141, 1027.1586, 1027.11, 1027.043, 1026.9829, 1026.919, 1026.8274, 1026.7389, 1026.6414, 1026.5344, 1026.4203, 1026.2593, 1026.1039, 1025.9264, 1025.7489, 1025.6506, 1025.4945, 1025.4106, 1025.2424, 1025.0964, 1024.972, 1024.8315, 1024.6174, 1024.5254, 1024.4417, 1024.3353, 1024.2524, 1024.2047, 1024.1395, 1024.0848, 1023.8707, 1023.7027, 1023.68506, NaN, NaN, 1029.2007, 1029.1719, 1029.1327, 1029.0851, 1029.0358, 1028.991, 1028.9424, 1028.8899, 1028.8436, 1028.7999, 1028.7562, 1028.709, 1028.6578, 1028.6115, 1028.5616, 1028.5117, 1028.4604, 1028.4098, 1028.365, 1028.3157, 1028.2648, 1028.2156, 1028.1678, 1028.1139, 1028.0623, 1028.012, 1027.9629, 1027.9075, 1027.8538, 1027.7985, 1027.7513, 1027.7015, 1027.6475, 1027.5925, 1027.5344, 1027.4697, 1027.4078, 1027.351, 1027.2963, 1027.2449, 1027.188, 1027.1362, 1027.0646, 1027.0, 1026.9224, 1026.8407, 1026.7363, 1026.6617, 1026.5889, 1026.48, 1026.3379, 1026.2257, 1026.1208, 1025.9897, 1025.8536, 1025.6846, 1025.5995, 1025.5015, 1025.3768, 1025.21, 1025.0668, 1024.9055, 1024.6208, 1024.5197, 1024.4856, 1024.4155, 1024.3153, 1024.2135, 1024.1217, 1023.866, 1023.68396, 1023.6627, NaN, NaN, 1029.2216, 1029.1921, 1029.1558, 1029.1019, 1029.0476, 1028.9916, 1028.9414, 1028.8922, 1028.8391, 1028.7874, 1028.7391, 1028.6866, 1028.634, 1028.5809, 1028.5303, 1028.4847, 1028.43, 1028.3806, 1028.3309, 1028.2751, 1028.2277, 1028.1732, 1028.1229, 1028.0725, 1028.0175, 1027.9587, 1027.8961, 1027.8463, 1027.7921, 1027.7437, 1027.6908, 1027.6414, 1027.5896, 1027.5431, 1027.4923, 1027.4446, 1027.3931, 1027.3414, 1027.2811, 1027.2163, 1027.1608, 1027.0931, 1027.0298, 1026.9602, 1026.8765, 1026.8079, 1026.7125, 1026.6041, 1026.4993, 1026.3861, 1026.2511, 1026.1461, 1025.9983, 1025.8112, 1025.717, 1025.6024, 1025.4369, 1025.3413, 1025.1649, 1024.9373, 1024.7709, 1024.5935, 1024.4415, 1024.3915, 1024.2938, 1024.2212, 1024.144, 1023.8099, 1023.6585, 1023.64026, NaN, NaN, 1029.2355, 1029.2091, 1029.1736, 1029.1194, 1029.0723, 1029.0212, 1028.9745, 1028.9235, 1028.8761, 1028.8284, 1028.7778, 1028.7238, 1028.6777, 1028.6261, 1028.5807, 1028.5394, 1028.497, 1028.4498, 1028.4088, 1028.363, 1028.3112, 1028.2546, 1028.1997, 1028.1523, 1028.1086, 1028.0642, 1028.0123, 1027.9539, 1027.9075, 1027.8589, 1027.8081, 1027.7615, 1027.7076, 1027.661, 1027.6147, 1027.5707, 1027.5138, 1027.4606, 1027.4082, 1027.3572, 1027.3007, 1027.2426, 1027.1826, 1027.1248, 1027.06, 1026.9974, 1026.9333, 1026.8767, 1026.8152, 1026.74, 1026.6558, 1026.577, 1026.4567, 1026.3247, 1026.1692, 1025.9893, 1025.7948, 1025.6501, 1025.534, 1025.3993, 1025.2856, 1025.1562, 1025.0083, 1024.7959, 1024.6324, 1024.5074, 1024.3827, 1024.3204, 1024.2454, 1024.1453, 1024.0343, 1023.6947, 1023.66266, 1023.64, 1023.6279, NaN, NaN, 1029.2029, 1029.1738, 1029.1351, 1029.0908, 1029.0422, 1028.9948, 1028.9487, 1028.8989, 1028.8525, 1028.8038, 1028.7548, 1028.703, 1028.656, 1028.6024, 1028.5454, 1028.4921, 1028.4408, 1028.39, 1028.3356, 1028.2808, 1028.2278, 1028.1742, 1028.1167, 1028.0624, 1028.0038, 1027.9478, 1027.8932, 1027.832, 1027.7731, 1027.729, 1027.6683, 1027.6152, 1027.5668, 1027.5049, 1027.4496, 1027.392, 1027.3239, 1027.2505, 1027.1968, 1027.1501, 1027.1056, 1027.0497, 1026.9778, 1026.8794, 1026.8104, 1026.752, 1026.6425, 1026.5363, 1026.4081, 1026.2607, 1026.0883, 1025.8618, 1025.6571, 1025.4979, 1025.409, 1025.3345, 1025.2374, 1025.1022, 1024.982, 1024.8575, 1024.6711, 1024.4921, 1024.3735, 1024.2574, 1024.1257, 1023.9116, 1023.7101, 1023.69073, 1023.6653, NaN, NaN, 1029.1959, 1029.166, 1029.1332, 1029.0878, 1029.0447, 1028.9968, 1028.9473, 1028.9043, 1028.8604, 1028.8147, 1028.769, 1028.7255, 1028.678, 1028.6327, 1028.5914, 1028.5404, 1028.4905, 1028.4414, 1028.3948, 1028.348, 1028.2955, 1028.2482, 1028.2007, 1028.1489, 1028.1023, 1028.0476, 1027.9958, 1027.9491, 1027.8987, 1027.8458, 1027.7938, 1027.7467, 1027.7015, 1027.6472, 1027.5953, 1027.5488, 1027.4988, 1027.4453, 1027.379, 1027.3347, 1027.2926, 1027.2389, 1027.1792, 1027.125, 1027.0732, 1027.0101, 1026.92, 1026.8435, 1026.7963, 1026.7374, 1026.6632, 1026.5461, 1026.429, 1026.2988, 1026.1616, 1026.0321, 1025.8594, 1025.7228, 1025.5751, 1025.4457, 1025.3057, 1025.1647, 1025.0249, 1024.8773, 1024.7021, 1024.4636, 1024.3168, 1024.2375, 1024.06, 1023.74896, 1023.7235, 1023.69763, 1023.6758, NaN, NaN, 1029.2106, 1029.1844, 1029.1483, 1029.1034, 1029.0599, 1029.0131, 1028.9679, 1028.9268, 1028.8782, 1028.8333, 1028.7894, 1028.7416, 1028.6895, 1028.6346, 1028.5873, 1028.5402, 1028.4948, 1028.4509, 1028.4043, 1028.3579, 1028.3103, 1028.2657, 1028.2207, 1028.1638, 1028.1195, 1028.0698, 1028.0115, 1027.9545, 1027.9026, 1027.8431, 1027.7946, 1027.7429, 1027.6987, 1027.6572, 1027.6085, 1027.553, 1027.5021, 1027.4509, 1027.4038, 1027.3579, 1027.3027, 1027.2439, 1027.174, 1027.1239, 1027.0592, 1026.9924, 1026.9352, 1026.8793, 1026.8201, 1026.7394, 1026.6498, 1026.5536, 1026.4357, 1026.3298, 1026.1882, 1025.9966, 1025.8196, 1025.6954, 1025.5773, 1025.4125, 1025.3105, 1025.2368, 1025.1444, 1025.0361, 1024.9357, 1024.7278, 1024.5498, 1024.4297, 1024.2261, 1024.0311, 1023.7688, 1023.73444, 1023.70715, 1023.68823, NaN, NaN, 1029.2288, 1029.203, 1029.1722, 1029.1295, 1029.081, 1029.0393, 1028.9972, 1028.9454, 1028.8989, 1028.8512, 1028.8042, 1028.7537, 1028.705, 1028.6588, 1028.6051, 1028.5442, 1028.4938, 1028.4412, 1028.3878, 1028.3383, 1028.2902, 1028.2386, 1028.1836, 1028.1298, 1028.0729, 1028.0184, 1027.96, 1027.9048, 1027.8535, 1027.7944, 1027.7349, 1027.6855, 1027.631, 1027.5835, 1027.5404, 1027.4861, 1027.4291, 1027.373, 1027.326, 1027.2769, 1027.2141, 1027.1512, 1027.0941, 1027.0455, 1026.9879, 1026.9142, 1026.8309, 1026.7134, 1026.6234, 1026.5386, 1026.4406, 1026.3196, 1026.1686, 1026.0292, 1025.8579, 1025.7225, 1025.6128, 1025.4752, 1025.3762, 1025.2632, 1025.1628, 1025.0748, 1024.8959, 1024.6176, 1024.385, 1024.2019, 1024.0353, 1023.78705, 1023.743, 1023.72534, 1023.7019, 1023.6906, NaN, NaN, 1029.2191, 1029.1917, 1029.1577, 1029.103, 1029.0497, 1028.9929, 1028.9368, 1028.8853, 1028.8403, 1028.7883, 1028.7365, 1028.6859, 1028.6339, 1028.5812, 1028.5292, 1028.4775, 1028.4247, 1028.3698, 1028.3224, 1028.2761, 1028.219, 1028.1641, 1028.1141, 1028.0626, 1028.0049, 1027.9491, 1027.8925, 1027.834, 1027.7831, 1027.7367, 1027.6875, 1027.6323, 1027.5802, 1027.5283, 1027.4767, 1027.4196, 1027.3488, 1027.2964, 1027.2389, 1027.1876, 1027.1394, 1027.0785, 1026.9889, 1026.8988, 1026.8157, 1026.7156, 1026.6592, 1026.568, 1026.4657, 1026.3302, 1026.2373, 1026.077, 1025.909, 1025.739, 1025.5958, 1025.3666, 1025.2229, 1025.118, 1024.9558, 1024.762, 1024.6193, 1024.5135, 1024.2532, 1024.0945, 1023.82526, 1023.78, 1023.7507, 1023.733, 1023.7138, NaN, NaN, 1029.207, 1029.1766, 1029.1367, 1029.079, 1029.0289, 1028.9775, 1028.928, 1028.8777, 1028.8219, 1028.7723, 1028.7255, 1028.6837, 1028.6364, 1028.5869, 1028.5356, 1028.4888, 1028.4305, 1028.3768, 1028.3279, 1028.274, 1028.2197, 1028.1705, 1028.1183, 1028.0664, 1028.0078, 1027.9464, 1027.8987, 1027.844, 1027.7975, 1027.7488, 1027.6912, 1027.6338, 1027.5875, 1027.5426, 1027.5013, 1027.4543, 1027.413, 1027.356, 1027.3036, 1027.2509, 1027.2009, 1027.1497, 1027.0873, 1027.001, 1026.9146, 1026.8287, 1026.733, 1026.6318, 1026.5411, 1026.4487, 1026.3417, 1026.207, 1026.0784, 1025.9169, 1025.741, 1025.6128, 1025.4299, 1025.2428, 1025.1091, 1024.9788, 1024.8945, 1024.6616, 1024.3788, 1024.2872, 1024.2206, 1023.99396, 1023.82, 1023.8003, 1023.7697, 1023.75555, NaN, NaN, 1029.2264, 1029.203, 1029.1686, 1029.1206, 1029.0734, 1029.024, 1028.9768, 1028.9303, 1028.8778, 1028.8265, 1028.7833, 1028.734, 1028.6804, 1028.6299, 1028.5791, 1028.5334, 1028.4828, 1028.4315, 1028.3875, 1028.3386, 1028.2858, 1028.2328, 1028.1777, 1028.1252, 1028.0659, 1028.0098, 1027.955, 1027.891, 1027.8348, 1027.7839, 1027.7285, 1027.6691, 1027.6138, 1027.5615, 1027.505, 1027.453, 1027.4026, 1027.3561, 1027.297, 1027.2506, 1027.197, 1027.1372, 1027.0723, 1027.0029, 1026.9177, 1026.8406, 1026.7483, 1026.6278, 1026.5516, 1026.4547, 1026.3217, 1026.1576, 1026.0295, 1025.8763, 1025.6902, 1025.5209, 1025.3838, 1025.2388, 1025.1326, 1025.0204, 1024.8911, 1024.7113, 1024.4318, 1024.2882, 1024.1965, 1023.9541, 1023.8856, 1023.8602, 1023.8429, 1023.82324, NaN, NaN, 1029.2216, 1029.1919, 1029.1558, 1029.1108, 1029.0652, 1029.0153, 1028.9679, 1028.9214, 1028.8698, 1028.8196, 1028.7634, 1028.7148, 1028.662, 1028.6127, 1028.5641, 1028.5121, 1028.4652, 1028.4225, 1028.3749, 1028.3243, 1028.2728, 1028.218, 1028.1665, 1028.1166, 1028.0717, 1028.0245, 1027.9717, 1027.9235, 1027.867, 1027.8164, 1027.7628, 1027.7078, 1027.6667, 1027.6166, 1027.5638, 1027.5188, 1027.4606, 1027.4052, 1027.3484, 1027.2915, 1027.2203, 1027.1718, 1027.1104, 1027.0461, 1026.9908, 1026.8993, 1026.8152, 1026.748, 1026.6508, 1026.5453, 1026.4044, 1026.2849, 1026.1659, 1026.0331, 1025.8887, 1025.7485, 1025.5463, 1025.3765, 1025.2351, 1025.1115, 1025.0332, 1024.9174, 1024.6594, 1024.4025, 1024.2594, 1024.0143, 1023.91797, 1023.899, 1023.8714, 1023.8495, NaN, NaN, 1029.197, 1029.166, 1029.1315, 1029.0825, 1029.0402, 1028.9985, 1028.9512, 1028.9084, 1028.8633, 1028.8175, 1028.7731, 1028.7363, 1028.6904, 1028.6525, 1028.6086, 1028.5612, 1028.5149, 1028.4714, 1028.4271, 1028.38, 1028.337, 1028.2893, 1028.2439, 1028.201, 1028.1561, 1028.1084, 1028.0619, 1028.0146, 1027.9711, 1027.9208, 1027.8774, 1027.8348, 1027.794, 1027.7527, 1027.7053, 1027.6576, 1027.606, 1027.5632, 1027.5184, 1027.4674, 1027.4253, 1027.3809, 1027.3367, 1027.276, 1027.222, 1027.1602, 1027.1124, 1027.051, 1026.997, 1026.9059, 1026.8182, 1026.74, 1026.6237, 1026.5089, 1026.3904, 1026.2915, 1026.1942, 1026.0847, 1025.9614, 1025.7897, 1025.6797, 1025.4967, 1025.362, 1025.2368, 1025.1339, 1025.0409, 1024.9048, 1024.6943, 1024.4425, 1024.2971, 1024.0671, 1023.92365, 1023.89514, 1023.8732, 1023.8465, NaN, NaN, 1029.2014, 1029.1742, 1029.1404, 1029.0978, 1029.0542, 1029.0103, 1028.9574, 1028.9113, 1028.8649, 1028.8127, 1028.761, 1028.7085, 1028.6548, 1028.6035, 1028.5488, 1028.4971, 1028.4437, 1028.3916, 1028.34, 1028.2897, 1028.2386, 1028.1936, 1028.1432, 1028.086, 1028.0293, 1027.9784, 1027.9303, 1027.876, 1027.8198, 1027.7632, 1027.7019, 1027.6486, 1027.6012, 1027.5573, 1027.5157, 1027.47, 1027.4219, 1027.3788, 1027.3298, 1027.269, 1027.2194, 1027.1516, 1027.0878, 1027.0264, 1026.9518, 1026.8574, 1026.7676, 1026.6592, 1026.5793, 1026.4822, 1026.3717, 1026.2513, 1026.1313, 1025.9727, 1025.7848, 1025.5955, 1025.4639, 1025.3348, 1025.2279, 1025.1298, 1024.9883, 1024.8384, 1024.5669, 1024.2825, 1023.97864, 1023.9357, 1023.9057, 1023.8905, 1023.86633, 1023.84033, 1023.82874, NaN, NaN, 1029.2057, 1029.1737, 1029.1366, 1029.0857, 1029.0349, 1028.9836, 1028.9333, 1028.876, 1028.8196, 1028.7614, 1028.7133, 1028.6608, 1028.6106, 1028.5626, 1028.5164, 1028.46, 1028.4122, 1028.3628, 1028.3145, 1028.2643, 1028.2177, 1028.1748, 1028.119, 1028.0762, 1028.0322, 1027.9827, 1027.9355, 1027.8815, 1027.8245, 1027.7695, 1027.7142, 1027.6619, 1027.6198, 1027.5731, 1027.5284, 1027.4749, 1027.4244, 1027.3732, 1027.3177, 1027.2573, 1027.2054, 1027.155, 1027.0979, 1027.0375, 1026.9397, 1026.817, 1026.7097, 1026.6123, 1026.5032, 1026.3676, 1026.2617, 1026.1503, 1026.0426, 1025.8579, 1025.6643, 1025.4933, 1025.3413, 1025.2518, 1025.161, 1025.0221, 1024.8502, 1024.6564, 1024.4059, 1024.0668, 1023.9577, 1023.9339, 1023.9025, 1023.87463, 1023.8632, NaN, NaN, 1029.2142, 1029.184, 1029.1477, 1029.1013, 1029.0553, 1029.0126, 1028.9656, 1028.9154, 1028.8678, 1028.8243, 1028.7755, 1028.7277, 1028.6769, 1028.6337, 1028.5864, 1028.5376, 1028.4875, 1028.441, 1028.3905, 1028.3474, 1028.3013, 1028.2576, 1028.2043, 1028.1599, 1028.113, 1028.065, 1028.0201, 1027.9689, 1027.9187, 1027.8718, 1027.8207, 1027.7761, 1027.7356, 1027.69, 1027.6426, 1027.5907, 1027.5417, 1027.4968, 1027.4464, 1027.3917, 1027.3322, 1027.2688, 1027.2, 1027.124, 1027.0527, 1026.9915, 1026.9186, 1026.8364, 1026.7732, 1026.6713, 1026.56, 1026.4261, 1026.2797, 1026.2001, 1026.0756, 1025.91, 1025.7542, 1025.6095, 1025.457, 1025.3217, 1025.2257, 1025.1449, 1025.0452, 1024.917, 1024.6797, 1024.349, 1024.0825, 1024.0334, 1024.0148, 1023.9839, 1023.9579, 1023.9506, NaN, NaN, 1029.1947, 1029.1692, 1029.1301, 1029.0846, 1029.0438, 1029.0054, 1028.9629, 1028.9136, 1028.8702, 1028.8276, 1028.786, 1028.7415, 1028.6919, 1028.651, 1028.6073, 1028.563, 1028.5173, 1028.4706, 1028.4263, 1028.3793, 1028.3247, 1028.2759, 1028.2277, 1028.1737, 1028.1213, 1028.0737, 1028.0189, 1027.9622, 1027.9143, 1027.8656, 1027.8154, 1027.7599, 1027.7068, 1027.659, 1027.6162, 1027.5709, 1027.5242, 1027.4788, 1027.4309, 1027.3862, 1027.3378, 1027.2837, 1027.2195, 1027.1311, 1027.0479, 1026.9774, 1026.9105, 1026.85, 1026.7355, 1026.6318, 1026.5367, 1026.3925, 1026.3085, 1026.2249, 1026.1191, 1026.0049, 1025.8422, 1025.7457, 1025.6226, 1025.4812, 1025.3279, 1025.2382, 1025.1455, 1025.0334, 1024.9283, 1024.7501, 1024.4578, 1024.2142, 1024.1208, 1024.0962, 1024.0691, 1024.049, 1024.0309, NaN, NaN, 1029.2021, 1029.1794, 1029.145, 1029.0974, 1029.0516, 1029.0118, 1028.9705, 1028.93, 1028.8905, 1028.845, 1028.791, 1028.7444, 1028.7018, 1028.6519, 1028.6046, 1028.5576, 1028.5154, 1028.4722, 1028.4209, 1028.3806, 1028.3286, 1028.2792, 1028.231, 1028.1826, 1028.1354, 1028.0878, 1028.0377, 1027.9875, 1027.9391, 1027.89, 1027.8381, 1027.7909, 1027.7296, 1027.6809, 1027.6306, 1027.5801, 1027.5195, 1027.4622, 1027.4069, 1027.3553, 1027.291, 1027.2332, 1027.1625, 1027.0957, 1027.0374, 1026.969, 1026.8921, 1026.8073, 1026.7139, 1026.6113, 1026.5023, 1026.3895, 1026.2819, 1026.196, 1026.0544, 1025.8883, 1025.7533, 1025.6628, 1025.4661, 1025.3308, 1025.2115, 1025.0969, 1024.9891, 1024.8601, 1024.6338, 1024.343, 1024.2377, 1024.2009, 1024.1732, 1024.1461, 1024.1207, 1024.1018, NaN, NaN, 1029.2113, 1029.1815, 1029.1396, 1029.0818, 1029.0282, 1028.9795, 1028.9335, 1028.8876, 1028.8408, 1028.7946, 1028.7428, 1028.6892, 1028.6302, 1028.5886, 1028.5371, 1028.4836, 1028.4305, 1028.3837, 1028.3354, 1028.2832, 1028.2365, 1028.1892, 1028.1389, 1028.0903, 1028.0392, 1027.9836, 1027.9337, 1027.8793, 1027.8236, 1027.7716, 1027.7137, 1027.654, 1027.5981, 1027.5497, 1027.4934, 1027.4335, 1027.3766, 1027.3228, 1027.259, 1027.1906, 1027.1155, 1027.0487, 1026.9982, 1026.9138, 1026.8143, 1026.6874, 1026.5848, 1026.5099, 1026.4255, 1026.3094, 1026.2029, 1026.0709, 1025.9098, 1025.7854, 1025.714, 1025.5385, 1025.3033, 1025.2175, 1025.1079, 1025.0112, 1024.9124, 1024.8273, 1024.5685, 1024.2544, 1024.2263, 1024.1976, 1024.182, 1024.1508, 1024.1261, NaN, NaN, 1029.2123, 1029.1895, 1029.1582, 1029.1111, 1029.0588, 1029.0096, 1028.9628, 1028.9144, 1028.8693, 1028.8192, 1028.7704, 1028.723, 1028.6741, 1028.6232, 1028.5714, 1028.5216, 1028.471, 1028.4246, 1028.3749, 1028.3219, 1028.272, 1028.224, 1028.1714, 1028.1233, 1028.0747, 1028.0273, 1027.9781, 1027.923, 1027.8713, 1027.8176, 1027.7533, 1027.69, 1027.6344, 1027.5735, 1027.5085, 1027.4503, 1027.3905, 1027.3375, 1027.2781, 1027.2258, 1027.16, 1027.0972, 1027.0272, 1026.9554, 1026.8856, 1026.7985, 1026.7, 1026.596, 1026.4884, 1026.3779, 1026.2556, 1026.1151, 1025.9967, 1025.7655, 1025.5596, 1025.3611, 1025.2544, 1025.1226, 1025.0314, 1024.9543, 1024.8295, 1024.4583, 1024.2639, 1024.2296, 1024.2036, 1024.1808, 1024.158, 1024.1385, 1024.1251, NaN, NaN, 1029.2112, 1029.1799, 1029.1449, 1029.0979, 1029.0543, 1029.0107, 1028.9685, 1028.9248, 1028.8741, 1028.8291, 1028.7817, 1028.7338, 1028.6846, 1028.6395, 1028.5918, 1028.5375, 1028.489, 1028.445, 1028.3917, 1028.3439, 1028.2924, 1028.2373, 1028.1943, 1028.1444, 1028.093, 1028.0466, 1027.9994, 1027.9563, 1027.9115, 1027.8674, 1027.8208, 1027.7734, 1027.7257, 1027.682, 1027.6318, 1027.5863, 1027.5359, 1027.4907, 1027.4344, 1027.3766, 1027.3254, 1027.2715, 1027.21, 1027.1451, 1027.0898, 1027.0098, 1026.9385, 1026.8612, 1026.7742, 1026.6538, 1026.5758, 1026.4908, 1026.3816, 1026.2522, 1026.1329, 1026.0116, 1025.8322, 1025.6691, 1025.5433, 1025.4536, 1025.3944, 1025.2908, 1025.2029, 1025.1133, 1025.0122, 1024.9023, 1024.7753, 1024.4902, 1024.2567, 1024.2076, 1024.17, 1024.1439, 1024.1296, 1024.1134, NaN, NaN, 1029.2117, 1029.1797, 1029.1427, 1029.0924, 1029.0469, 1029.0021, 1028.955, 1028.9052, 1028.8566, 1028.8088, 1028.76, 1028.7091, 1028.6646, 1028.6213, 1028.5762, 1028.5256, 1028.4797, 1028.4362, 1028.3942, 1028.3436, 1028.2932, 1028.2429, 1028.2006, 1028.1497, 1028.101, 1028.0537, 1028.0074, 1027.9633, 1027.9135, 1027.8597, 1027.8141, 1027.7671, 1027.7131, 1027.6628, 1027.6102, 1027.5613, 1027.5073, 1027.4493, 1027.3905, 1027.3367, 1027.2828, 1027.2236, 1027.162, 1027.0936, 1027.0297, 1026.9742, 1026.9099, 1026.8379, 1026.7584, 1026.68, 1026.5828, 1026.4952, 1026.3788, 1026.283, 1026.1823, 1026.0576, 1025.8794, 1025.6946, 1025.5613, 1025.416, 1025.3025, 1025.1843, 1025.1135, 1025.023, 1024.9266, 1024.7957, 1024.3734, 1024.2451, 1024.202, 1024.182, 1024.1592, 1024.1367, NaN, NaN, 1029.203, 1029.1726, 1029.136, 1029.0885, 1029.0339, 1028.981, 1028.9308, 1028.8826, 1028.8341, 1028.7853, 1028.7356, 1028.6826, 1028.6268, 1028.5768, 1028.528, 1028.4803, 1028.4323, 1028.3855, 1028.3379, 1028.2883, 1028.2385, 1028.1953, 1028.1447, 1028.0948, 1028.0457, 1027.9965, 1027.9475, 1027.9008, 1027.8492, 1027.8, 1027.7483, 1027.6919, 1027.6305, 1027.5726, 1027.5205, 1027.4646, 1027.397, 1027.3405, 1027.2875, 1027.2225, 1027.1549, 1027.0936, 1027.0314, 1026.9609, 1026.8901, 1026.8075, 1026.7526, 1026.6807, 1026.5946, 1026.5107, 1026.4044, 1026.2981, 1026.1863, 1026.0674, 1025.9136, 1025.7428, 1025.5494, 1025.4006, 1025.2457, 1025.1239, 1024.9825, 1024.7488, 1024.3885, 1024.3029, 1024.26, 1024.2351, 1024.2153, 1024.1823, 1024.164, 1024.1483, NaN, NaN, 1029.2115, 1029.1875, 1029.15, 1029.1, 1029.0499, 1029.0002, 1028.9486, 1028.8966, 1028.8431, 1028.7919, 1028.7439, 1028.6873, 1028.6362, 1028.5903, 1028.5457, 1028.4998, 1028.4539, 1028.4033, 1028.3527, 1028.3033, 1028.2573, 1028.2142, 1028.1666, 1028.114, 1028.0659, 1028.019, 1027.9677, 1027.9211, 1027.8755, 1027.8214, 1027.7723, 1027.7288, 1027.6835, 1027.6439, 1027.597, 1027.5428, 1027.4911, 1027.4425, 1027.3857, 1027.3391, 1027.2904, 1027.2418, 1027.1826, 1027.1174, 1027.0526, 1026.9774, 1026.9001, 1026.8185, 1026.737, 1026.6396, 1026.5426, 1026.4336, 1026.2782, 1026.1152, 1025.9424, 1025.776, 1025.6373, 1025.5658, 1025.4723, 1025.271, 1025.1536, 1025.085, 1025.0032, 1024.8682, 1024.5363, 1024.3657, 1024.3236, 1024.2865, 1024.2582, 1024.2329, 1024.2086, 1024.1901, NaN, NaN, 1029.235, 1029.2092, 1029.1703, 1029.1189, 1029.0685, 1029.0166, 1028.9635, 1028.9131, 1028.8615, 1028.809, 1028.7568, 1028.7053, 1028.6504, 1028.5979, 1028.5468, 1028.4957, 1028.4479, 1028.396, 1028.35, 1028.3007, 1028.2509, 1028.2079, 1028.1573, 1028.1019, 1028.046, 1027.9958, 1027.9503, 1027.9052, 1027.856, 1027.8036, 1027.7533, 1027.7054, 1027.6593, 1027.5978, 1027.5475, 1027.495, 1027.4347, 1027.3833, 1027.325, 1027.2549, 1027.1678, 1027.098, 1027.0453, 1026.9966, 1026.9375, 1026.8768, 1026.8193, 1026.7327, 1026.6733, 1026.6082, 1026.5317, 1026.3983, 1026.2181, 1026.0813, 1025.9415, 1025.7689, 1025.6241, 1025.4685, 1025.2577, 1025.1002, 1025.0033, 1024.8789, 1024.5417, 1024.3712, 1024.3468, 1024.3219, 1024.2942, 1024.2715, 1024.2511, 1024.2336, 1024.2201, NaN, NaN, 1029.2098, 1029.1846, 1029.1477, 1029.104, 1029.0604, 1029.0137, 1028.9681, 1028.9205, 1028.8745, 1028.8247, 1028.776, 1028.7314, 1028.6875, 1028.6417, 1028.593, 1028.5447, 1028.4943, 1028.4502, 1028.4033, 1028.361, 1028.3173, 1028.2704, 1028.2269, 1028.1733, 1028.1218, 1028.0693, 1028.0134, 1027.9633, 1027.9122, 1027.8566, 1027.8085, 1027.7631, 1027.712, 1027.6492, 1027.5961, 1027.547, 1027.4882, 1027.4348, 1027.3877, 1027.3322, 1027.2616, 1027.189, 1027.141, 1027.0748, 1027.0017, 1026.9333, 1026.8807, 1026.8075, 1026.7273, 1026.6655, 1026.5753, 1026.4507, 1026.351, 1026.2648, 1026.1332, 1026.0449, 1025.9006, 1025.729, 1025.593, 1025.4497, 1025.311, 1025.1305, 1024.9833, 1024.8353, 1024.508, 1024.3508, 1024.3243, 1024.3021, 1024.2786, 1024.2507, 1024.2325, NaN, NaN, 1029.2078, 1029.1788, 1029.144, 1029.0908, 1029.0365, 1028.9862, 1028.9352, 1028.8768, 1028.8218, 1028.7745, 1028.7291, 1028.678, 1028.6282, 1028.582, 1028.5271, 1028.4786, 1028.4385, 1028.3923, 1028.347, 1028.3063, 1028.2573, 1028.2057, 1028.1586, 1028.0981, 1028.0424, 1027.9941, 1027.9447, 1027.8832, 1027.834, 1027.7832, 1027.7329, 1027.6738, 1027.6249, 1027.5762, 1027.5354, 1027.4764, 1027.4235, 1027.3684, 1027.3058, 1027.2457, 1027.1772, 1027.1038, 1027.0166, 1026.94, 1026.8466, 1026.7678, 1026.6844, 1026.5917, 1026.4962, 1026.3749, 1026.266, 1026.1404, 1026.0103, 1025.8861, 1025.7051, 1025.5497, 1025.442, 1025.3247, 1025.2242, 1025.1167, 1025.0334, 1024.9286, 1024.7504, 1024.4307, 1024.3408, 1024.3146, 1024.2948, 1024.273, 1024.2533, 1024.2405, NaN, NaN, 1029.2081, 1029.1848, 1029.1539, 1029.1122, 1029.0721, 1029.0227, 1028.9786, 1028.9294, 1028.8784, 1028.8265, 1028.7795, 1028.727, 1028.6753, 1028.6288, 1028.5886, 1028.5466, 1028.5038, 1028.4589, 1028.4178, 1028.373, 1028.3236, 1028.2828, 1028.2399, 1028.1974, 1028.1538, 1028.1094, 1028.0607, 1028.0071, 1027.96, 1027.9169, 1027.8707, 1027.8264, 1027.7764, 1027.7263, 1027.675, 1027.6195, 1027.5653, 1027.5093, 1027.4545, 1027.3948, 1027.3295, 1027.2599, 1027.1921, 1027.1305, 1027.0629, 1026.99, 1026.9131, 1026.8303, 1026.7253, 1026.6486, 1026.537, 1026.406, 1026.3074, 1026.1985, 1026.0643, 1025.9021, 1025.7076, 1025.6106, 1025.4993, 1025.3905, 1025.2784, 1025.1649, 1025.0768, 1024.9823, 1024.8745, 1024.6681, 1024.3639, 1024.3235, 1024.301, 1024.2756, 1024.2493, 1024.2292, NaN, NaN, 1029.2308, 1029.205, 1029.1722, 1029.116, 1029.0667, 1029.017, 1028.9729, 1028.9235, 1028.8735, 1028.8188, 1028.7711, 1028.7188, 1028.6599, 1028.6046, 1028.5514, 1028.4999, 1028.4491, 1028.4009, 1028.3527, 1028.3027, 1028.2474, 1028.1957, 1028.1477, 1028.0917, 1028.0393, 1027.988, 1027.9355, 1027.8822, 1027.8325, 1027.7786, 1027.7313, 1027.6763, 1027.6217, 1027.5662, 1027.5088, 1027.4535, 1027.3865, 1027.3247, 1027.2732, 1027.2137, 1027.1522, 1027.0779, 1027.0051, 1026.9335, 1026.863, 1026.789, 1026.6813, 1026.5687, 1026.4905, 1026.3812, 1026.2811, 1026.1158, 1025.9539, 1025.7822, 1025.6292, 1025.4902, 1025.353, 1025.298, 1025.203, 1025.0771, 1024.9576, 1024.8223, 1024.6768, 1024.3666, 1024.3196, 1024.2921, 1024.2605, 1024.2281, NaN, NaN, 1029.2365, 1029.21, 1029.1707, 1029.1168, 1029.0631, 1029.014, 1028.9657, 1028.9193, 1028.8733, 1028.8293, 1028.7883, 1028.7362, 1028.6874, 1028.645, 1028.5958, 1028.5504, 1028.5024, 1028.4554, 1028.4043, 1028.3529, 1028.2981, 1028.2477, 1028.1968, 1028.1484, 1028.0964, 1028.041, 1027.9841, 1027.9287, 1027.8782, 1027.8313, 1027.776, 1027.7295, 1027.6727, 1027.6241, 1027.5691, 1027.512, 1027.449, 1027.3868, 1027.3246, 1027.2614, 1027.1957, 1027.137, 1027.0745, 1027.0004, 1026.9386, 1026.8523, 1026.7649, 1026.657, 1026.5308, 1026.4117, 1026.2958, 1026.1678, 1026.0916, 1025.9205, 1025.7651, 1025.6445, 1025.5426, 1025.4381, 1025.3429, 1025.2336, 1025.1339, 1025.0403, 1024.8986, 1024.7487, 1024.4252, 1024.3601, 1024.3385, 1024.3143, 1024.29, 1024.2559, 1024.2156, 1024.1753, NaN, NaN, 1029.206, 1029.178, 1029.145, 1029.0977, 1029.0555, 1029.006, 1028.9592, 1028.9081, 1028.8523, 1028.7983, 1028.7504, 1028.7079, 1028.6628, 1028.6088, 1028.5631, 1028.514, 1028.4642, 1028.4163, 1028.3677, 1028.3197, 1028.2703, 1028.2168, 1028.1664, 1028.119, 1028.0688, 1028.0176, 1027.9717, 1027.915, 1027.8622, 1027.8055, 1027.7495, 1027.6956, 1027.6486, 1027.5946, 1027.5426, 1027.4927, 1027.441, 1027.3745, 1027.3115, 1027.2499, 1027.1868, 1027.1089, 1027.047, 1026.979, 1026.9075, 1026.7822, 1026.6998, 1026.582, 1026.4489, 1026.3438, 1026.1903, 1026.0166, 1025.8904, 1025.7694, 1025.6011, 1025.46, 1025.3231, 1025.2128, 1025.1056, 1025.0216, 1024.8827, 1024.6979, 1024.3696, 1024.3137, 1024.2877, 1024.2592, 1024.2174, 1024.1561, 1024.1381, NaN, NaN, 1029.1967, 1029.173, 1029.1393, 1029.0895, 1029.0447, 1028.9988, 1028.9552, 1028.9071, 1028.8595, 1028.8108, 1028.7631, 1028.7173, 1028.6705, 1028.6229, 1028.5739, 1028.5187, 1028.4692, 1028.4235, 1028.3767, 1028.3256, 1028.272, 1028.2216, 1028.1708, 1028.1288, 1028.0837, 1028.0342, 1027.9819, 1027.9387, 1027.8928, 1027.8463, 1027.8018, 1027.752, 1027.6981, 1027.6459, 1027.5969, 1027.551, 1027.4929, 1027.4344, 1027.3812, 1027.3304, 1027.2709, 1027.2162, 1027.1371, 1027.0724, 1026.967, 1026.8801, 1026.8018, 1026.7462, 1026.6816, 1026.57, 1026.4202, 1026.3175, 1026.2163, 1026.1113, 1025.973, 1025.8086, 1025.7013, 1025.5613, 1025.4319, 1025.3207, 1025.2515, 1025.115, 1025.0088, 1024.9044, 1024.7509, 1024.5044, 1024.2615, 1024.2375, 1024.2113, 1024.1853, 1024.1428, 1024.0745, 1024.0375, NaN, NaN, 1029.2003, 1029.1732, 1029.1376, 1029.0944, 1029.046, 1028.9968, 1028.9512, 1028.9028, 1028.8557, 1028.8091, 1028.7627, 1028.717, 1028.6722, 1028.6227, 1028.5748, 1028.53, 1028.4777, 1028.4219, 1028.3723, 1028.3236, 1028.2728, 1028.2229, 1028.1702, 1028.1182, 1028.0708, 1028.0251, 1027.9757, 1027.9268, 1027.8793, 1027.8308, 1027.7802, 1027.727, 1027.6803, 1027.6295, 1027.5746, 1027.5138, 1027.4497, 1027.3947, 1027.3333, 1027.2793, 1027.2118, 1027.151, 1027.0751, 1027.0023, 1026.9346, 1026.8679, 1026.7865, 1026.7113, 1026.6486, 1026.5715, 1026.4843, 1026.3479, 1026.2278, 1026.059, 1025.9508, 1025.8164, 1025.6904, 1025.5585, 1025.4419, 1025.3036, 1025.1469, 1025.0264, 1024.8706, 1024.701, 1024.4283, 1024.19, 1024.1575, 1024.1293, 1024.1075, 1024.0793, 1024.0298, 1024.0049, NaN, NaN, 1029.2239, 1029.1981, 1029.1626, 1029.1127, 1029.057, 1029.0094, 1028.9565, 1028.9059, 1028.8495, 1028.7937, 1028.7375, 1028.686, 1028.6323, 1028.5834, 1028.5349, 1028.4835, 1028.4296, 1028.381, 1028.3304, 1028.2737, 1028.2156, 1028.1658, 1028.1182, 1028.0593, 1027.9984, 1027.9468, 1027.895, 1027.8406, 1027.7812, 1027.724, 1027.6674, 1027.6174, 1027.5603, 1027.5077, 1027.4526, 1027.4008, 1027.3484, 1027.2844, 1027.2323, 1027.1763, 1027.114, 1027.0433, 1026.972, 1026.8954, 1026.8147, 1026.7393, 1026.6675, 1026.5742, 1026.4803, 1026.3358, 1026.1903, 1026.0654, 1025.9359, 1025.7357, 1025.6053, 1025.4711, 1025.3469, 1025.2422, 1025.1327, 1025.0237, 1024.8918, 1024.6976, 1024.2958, 1024.1625, 1024.1309, 1024.0875, 1024.0396, 1024.0122, NaN, NaN, 1029.2075, 1029.1765, 1029.1398, 1029.089, 1029.0388, 1028.993, 1028.9458, 1028.8993, 1028.854, 1028.8116, 1028.759, 1028.7102, 1028.6646, 1028.6184, 1028.5771, 1028.5325, 1028.4857, 1028.4401, 1028.3898, 1028.3403, 1028.2921, 1028.2346, 1028.1769, 1028.1256, 1028.0774, 1028.0232, 1027.967, 1027.9056, 1027.847, 1027.7897, 1027.7314, 1027.6794, 1027.6252, 1027.5762, 1027.5226, 1027.4602, 1027.4039, 1027.3461, 1027.2902, 1027.2458, 1027.1959, 1027.1201, 1027.065, 1027.0071, 1026.9414, 1026.876, 1026.8038, 1026.7153, 1026.634, 1026.5314, 1026.4387, 1026.3438, 1026.2092, 1026.0765, 1025.9769, 1025.8428, 1025.724, 1025.5363, 1025.371, 1025.2448, 1025.1528, 1025.0286, 1024.9017, 1024.6703, 1024.2385, 1024.1527, 1024.1063, 1024.0548, 1024.0052, 1023.86096, 1023.8347, NaN, NaN, 1029.1995, 1029.1755, 1029.1476, 1029.0981, 1029.0522, 1029.0084, 1028.9663, 1028.9233, 1028.8777, 1028.8356, 1028.7833, 1028.7323, 1028.6859, 1028.6404, 1028.5889, 1028.534, 1028.4872, 1028.44, 1028.391, 1028.3362, 1028.2804, 1028.2234, 1028.1731, 1028.1182, 1028.0704, 1028.0223, 1027.9718, 1027.9226, 1027.8716, 1027.8179, 1027.7655, 1027.7156, 1027.6597, 1027.6038, 1027.545, 1027.4883, 1027.4365, 1027.3855, 1027.334, 1027.286, 1027.2316, 1027.1731, 1027.1012, 1027.041, 1026.9694, 1026.8871, 1026.794, 1026.7008, 1026.6162, 1026.5292, 1026.4072, 1026.2373, 1026.1172, 1026.0131, 1025.8503, 1025.7234, 1025.5846, 1025.4044, 1025.2677, 1025.1245, 1024.9996, 1024.8115, 1024.6654, 1024.2666, 1024.1208, 1024.0182, 1023.9385, 1023.85345, 1023.8091, 1023.79083, NaN, NaN, 1029.1774, 1029.1512, 1029.1145, 1029.0629, 1029.0162, 1028.9681, 1028.921, 1028.8782, 1028.8348, 1028.7891, 1028.737, 1028.6887, 1028.6401, 1028.589, 1028.5372, 1028.4895, 1028.4344, 1028.3829, 1028.3313, 1028.2784, 1028.2308, 1028.1772, 1028.125, 1028.0751, 1028.0168, 1027.964, 1027.9104, 1027.8595, 1027.8097, 1027.7565, 1027.7048, 1027.6522, 1027.5892, 1027.5377, 1027.4835, 1027.424, 1027.3619, 1027.3167, 1027.266, 1027.2036, 1027.1443, 1027.0576, 1026.9763, 1026.9193, 1026.859, 1026.7944, 1026.7097, 1026.6195, 1026.5046, 1026.3932, 1026.2761, 1026.1628, 1026.074, 1025.9203, 1025.723, 1025.6029, 1025.4902, 1025.4008, 1025.2928, 1025.1495, 1025.0289, 1024.9459, 1024.8597, 1024.6244, 1024.2025, 1024.0309, 1023.88196, 1023.81616, 1023.7845, 1023.75854, 1023.73755, NaN, NaN, 1029.2032, 1029.1791, 1029.1447, 1029.0939, 1029.0448, 1028.9941, 1028.9398, 1028.8867, 1028.8335, 1028.7842, 1028.7313, 1028.6831, 1028.6274, 1028.5737, 1028.5249, 1028.4695, 1028.4172, 1028.3644, 1028.3121, 1028.2615, 1028.2024, 1028.149, 1028.1011, 1028.0525, 1028.0055, 1027.9487, 1027.8987, 1027.8457, 1027.7935, 1027.7365, 1027.6835, 1027.6377, 1027.5829, 1027.5321, 1027.4764, 1027.4259, 1027.3644, 1027.2992, 1027.2416, 1027.1833, 1027.1158, 1027.0591, 1026.994, 1026.9325, 1026.8735, 1026.7855, 1026.7062, 1026.6373, 1026.556, 1026.4629, 1026.3524, 1026.2003, 1026.0195, 1025.9055, 1025.8058, 1025.6416, 1025.4841, 1025.3093, 1025.1833, 1025.0472, 1024.9102, 1024.7631, 1024.5165, 1024.0029, 1023.8356, 1023.7774, 1023.7383, 1023.7115, 1023.689, NaN, NaN, 1029.1965, 1029.1652, 1029.1343, 1029.0902, 1029.0438, 1029.0009, 1028.956, 1028.9147, 1028.8683, 1028.8207, 1028.772, 1028.7255, 1028.6781, 1028.6337, 1028.5884, 1028.543, 1028.5016, 1028.4564, 1028.4102, 1028.3674, 1028.3188, 1028.2748, 1028.2277, 1028.1833, 1028.1449, 1028.0894, 1028.0383, 1027.9907, 1027.932, 1027.8795, 1027.8248, 1027.7739, 1027.7158, 1027.6631, 1027.6104, 1027.5569, 1027.4989, 1027.4493, 1027.3972, 1027.337, 1027.2788, 1027.2238, 1027.1663, 1027.1102, 1027.0327, 1026.9606, 1026.8918, 1026.8163, 1026.731, 1026.6562, 1026.5542, 1026.4711, 1026.3855, 1026.2826, 1026.1791, 1026.073, 1025.9187, 1025.7837, 1025.6477, 1025.4819, 1025.2924, 1025.1342, 1025.0454, 1024.8752, 1024.5885, 1023.9839, 1023.92755, 1023.8686, 1023.73175, 1023.68665, 1023.6682, NaN, NaN, 1029.1768, 1029.1472, 1029.11, 1029.0674, 1029.029, 1028.9816, 1028.9358, 1028.891, 1028.8383, 1028.7948, 1028.7539, 1028.7078, 1028.6594, 1028.6215, 1028.575, 1028.5292, 1028.4802, 1028.4354, 1028.3892, 1028.345, 1028.295, 1028.2375, 1028.1858, 1028.137, 1028.0944, 1028.0474, 1027.9836, 1027.9354, 1027.8909, 1027.853, 1027.7927, 1027.7434, 1027.6974, 1027.6548, 1027.6062, 1027.5516, 1027.5046, 1027.442, 1027.3804, 1027.3214, 1027.2659, 1027.2012, 1027.1473, 1027.0969, 1027.0442, 1026.9933, 1026.9451, 1026.8948, 1026.8358, 1026.7856, 1026.7366, 1026.6794, 1026.6122, 1026.5247, 1026.4124, 1026.3085, 1026.2043, 1026.0724, 1025.98, 1025.8777, 1025.7007, 1025.5447, 1025.3824, 1025.2198, 1025.0786, 1024.904, 1024.6674, 1024.3427, 1023.95483, 1023.90497, 1023.76746, 1023.6983, 1023.675, 1023.65924, NaN, NaN, 1029.1893, 1029.1661, 1029.1327, 1029.0881, 1029.0356, 1028.9874, 1028.9362, 1028.8829, 1028.8303, 1028.7765, 1028.7246, 1028.6678, 1028.6139, 1028.5635, 1028.5093, 1028.449, 1028.3981, 1028.3469, 1028.2942, 1028.2426, 1028.1849, 1028.1388, 1028.0865, 1028.0319, 1027.9836, 1027.9335, 1027.8812, 1027.8258, 1027.7611, 1027.7054, 1027.6515, 1027.5974, 1027.5283, 1027.4708, 1027.4001, 1027.3374, 1027.27, 1027.2172, 1027.168, 1027.1095, 1027.0531, 1026.993, 1026.9333, 1026.8737, 1026.8073, 1026.738, 1026.6559, 1026.5691, 1026.4614, 1026.3348, 1026.2158, 1026.0898, 1025.9629, 1025.8062, 1025.6437, 1025.5233, 1025.3167, 1025.1431, 1024.9783, 1024.762, 1024.1777, 1023.95966, 1023.9212, 1023.8492, 1023.7486, 1023.7222, 1023.697, 1023.6836, NaN, NaN, 1029.1449, 1029.1174, 1029.0844, 1029.0408, 1028.9954, 1028.9469, 1028.9009, 1028.8518, 1028.8036, 1028.7528, 1028.7072, 1028.657, 1028.6027, 1028.552, 1028.5073, 1028.4628, 1028.4146, 1028.3687, 1028.3157, 1028.2599, 1028.2085, 1028.1542, 1028.093, 1028.0371, 1027.9766, 1027.9298, 1027.8705, 1027.8234, 1027.7687, 1027.6986, 1027.6257, 1027.5532, 1027.4835, 1027.4146, 1027.354, 1027.2991, 1027.2365, 1027.1774, 1027.1206, 1027.0641, 1027.0126, 1026.962, 1026.9087, 1026.8528, 1026.7919, 1026.7283, 1026.6659, 1026.5944, 1026.505, 1026.4114, 1026.3096, 1026.1584, 1025.9773, 1025.8185, 1025.627, 1025.4396, 1025.2853, 1025.0785, 1024.8256, 1024.6477, 1024.1144, 1023.9307, 1023.90643, 1023.82007, 1023.73346, 1023.70667, NaN, NaN, 1029.1693, 1029.1423, 1029.1083, 1029.0658, 1029.0225, 1028.9823, 1028.937, 1028.8947, 1028.8549, 1028.8142, 1028.7725, 1028.7305, 1028.6838, 1028.6407, 1028.5972, 1028.557, 1028.5162, 1028.4681, 1028.4263, 1028.381, 1028.3342, 1028.2819, 1028.2296, 1028.181, 1028.124, 1028.0791, 1028.0261, 1027.978, 1027.9237, 1027.8514, 1027.7761, 1027.7166, 1027.6538, 1027.5906, 1027.5269, 1027.4716, 1027.4043, 1027.3342, 1027.268, 1027.2135, 1027.1669, 1027.121, 1027.0763, 1027.0299, 1026.9818, 1026.935, 1026.8933, 1026.8518, 1026.8077, 1026.7563, 1026.7054, 1026.6365, 1026.531, 1026.379, 1026.2607, 1026.1322, 1025.9585, 1025.8223, 1025.6978, 1025.5482, 1025.3853, 1025.2366, 1025.0569, 1024.9307, 1024.6945, 1024.2318, 1023.84033, 1023.8069, 1023.78937, 1023.7706, 1023.75653, NaN, NaN, 1029.1819, 1029.1617, 1029.133, 1029.0876, 1029.0454, 1029.0015, 1028.9523, 1028.904, 1028.8563, 1028.8069, 1028.7557, 1028.7024, 1028.6552, 1028.6077, 1028.5643, 1028.5205, 1028.4764, 1028.4296, 1028.3839, 1028.339, 1028.2986, 1028.2554, 1028.2129, 1028.1694, 1028.1223, 1028.0721, 1028.0198, 1027.966, 1027.9175, 1027.8601, 1027.7954, 1027.741, 1027.6622, 1027.6013, 1027.5413, 1027.4825, 1027.417, 1027.359, 1027.3003, 1027.2437, 1027.1882, 1027.1357, 1027.083, 1027.0267, 1026.9773, 1026.9252, 1026.8824, 1026.8383, 1026.7954, 1026.7476, 1026.7059, 1026.6487, 1026.5629, 1026.4891, 1026.3912, 1026.2034, 1026.0787, 1025.9242, 1025.6993, 1025.5096, 1025.4005, 1025.2732, 1025.1418, 1025.0288, 1024.9225, 1024.7257, 1024.2742, 1023.8938, 1023.8605, 1023.8371, 1023.81134, 1023.79144, 1023.7784, NaN, NaN, 1029.1752, 1029.1525, 1029.1189, 1029.0685, 1029.0239, 1028.9752, 1028.9264, 1028.8806, 1028.8259, 1028.7728, 1028.7233, 1028.6758, 1028.6241, 1028.5829, 1028.5413, 1028.4911, 1028.4426, 1028.3966, 1028.3549, 1028.3047, 1028.2571, 1028.2058, 1028.1575, 1028.0988, 1028.0465, 1027.9993, 1027.9557, 1027.9016, 1027.8451, 1027.7571, 1027.6686, 1027.6152, 1027.5494, 1027.4937, 1027.4369, 1027.3696, 1027.3148, 1027.2501, 1027.1985, 1027.1552, 1027.1124, 1027.0668, 1027.0197, 1026.9695, 1026.9263, 1026.8821, 1026.8339, 1026.7837, 1026.7406, 1026.682, 1026.6057, 1026.5536, 1026.4762, 1026.3347, 1026.1471, 1026.0027, 1025.8702, 1025.7379, 1025.5844, 1025.4523, 1025.2869, 1025.1165, 1024.9789, 1024.8416, 1024.6923, 1024.4222, 1023.87, 1023.8166, 1023.79834, 1023.78094, NaN, NaN, 1029.1775, 1029.1499, 1029.1128, 1029.0718, 1029.0323, 1028.9884, 1028.9478, 1028.9034, 1028.8544, 1028.8021, 1028.7557, 1028.7096, 1028.6616, 1028.6147, 1028.5675, 1028.5231, 1028.4805, 1028.4348, 1028.3871, 1028.3389, 1028.288, 1028.2363, 1028.1788, 1028.1254, 1028.0734, 1028.0096, 1027.957, 1027.911, 1027.8457, 1027.7722, 1027.6919, 1027.623, 1027.5605, 1027.5009, 1027.4398, 1027.3732, 1027.3094, 1027.2552, 1027.1976, 1027.1547, 1027.1093, 1027.0566, 1027.0162, 1026.9702, 1026.93, 1026.8907, 1026.8444, 1026.8003, 1026.7554, 1026.7113, 1026.6584, 1026.601, 1026.5504, 1026.4749, 1026.3341, 1026.1952, 1025.9282, 1025.6484, 1025.3617, 1025.2247, 1025.1201, 1024.9559, 1024.7703, 1024.4979, 1024.0325, 1023.8444, 1023.8188, 1023.799, 1023.77527, 1023.75226, NaN, NaN, 1029.1617, 1029.1365, 1029.1028, 1029.0586, 1029.0181, 1028.974, 1028.929, 1028.884, 1028.8425, 1028.8002, 1028.7599, 1028.7188, 1028.6786, 1028.6388, 1028.6001, 1028.5574, 1028.5133, 1028.4714, 1028.4313, 1028.3923, 1028.354, 1028.2988, 1028.256, 1028.2169, 1028.1658, 1028.1157, 1028.0657, 1028.017, 1027.953, 1027.8865, 1027.8326, 1027.7833, 1027.727, 1027.6587, 1027.6119, 1027.5563, 1027.4795, 1027.4342, 1027.3752, 1027.3153, 1027.2511, 1027.2054, 1027.1593, 1027.1139, 1027.0673, 1027.016, 1026.9733, 1026.931, 1026.8862, 1026.84, 1026.7977, 1026.7543, 1026.7041, 1026.6384, 1026.583, 1026.5308, 1026.4528, 1026.3242, 1026.21, 1026.0482, 1025.8679, 1025.706, 1025.5022, 1025.3304, 1025.2512, 1025.0739, 1024.9476, 1024.8011, 1024.5515, 1023.9599, 1023.8502, 1023.81744, 1023.7902, 1023.76044, 1023.7426, NaN, NaN, 1029.1879, 1029.1647, 1029.1323, 1029.0875, 1029.0377, 1028.9907, 1028.9425, 1028.8962, 1028.8478, 1028.8005, 1028.7505, 1028.7025, 1028.6516, 1028.6001, 1028.5482, 1028.4973, 1028.4432, 1028.3904, 1028.3402, 1028.2863, 1028.2306, 1028.1754, 1028.1215, 1028.0574, 1027.998, 1027.9293, 1027.8739, 1027.8214, 1027.7616, 1027.7058, 1027.6492, 1027.5917, 1027.5255, 1027.4587, 1027.4067, 1027.3495, 1027.2897, 1027.2268, 1027.1658, 1027.1094, 1027.0531, 1027.0012, 1026.9506, 1026.8995, 1026.8462, 1026.7914, 1026.7347, 1026.6669, 1026.5875, 1026.514, 1026.4148, 1026.2877, 1026.1779, 1026.0652, 1025.8955, 1025.6665, 1025.4346, 1025.2947, 1025.1696, 1025.0638, 1024.9652, 1024.8104, 1024.301, 1023.8869, 1023.8336, 1023.80756, 1023.7785, 1023.7448, 1023.72424, NaN, NaN, 1029.1841, 1029.1588, 1029.1267, 1029.0787, 1029.0332, 1028.9895, 1028.9425, 1028.8928, 1028.8478, 1028.803, 1028.7562, 1028.7101, 1028.6655, 1028.6256, 1028.5778, 1028.5316, 1028.4857, 1028.4419, 1028.3878, 1028.3422, 1028.2963, 1028.2439, 1028.1965, 1028.1394, 1028.0911, 1028.0436, 1027.9861, 1027.9294, 1027.8785, 1027.8252, 1027.759, 1027.7057, 1027.659, 1027.6067, 1027.5558, 1027.4895, 1027.4194, 1027.3552, 1027.2883, 1027.2379, 1027.1859, 1027.136, 1027.084, 1027.0273, 1026.9738, 1026.9269, 1026.8688, 1026.8059, 1026.7458, 1026.6752, 1026.6011, 1026.519, 1026.4285, 1026.2883, 1026.1705, 1026.0316, 1025.9088, 1025.7871, 1025.6631, 1025.4664, 1025.2896, 1025.1617, 1025.0468, 1024.9181, 1024.7288, 1024.2073, 1023.95044, 1023.9096, 1023.84875, 1023.7915, 1023.76605, 1023.7533, NaN, NaN, 1029.1852, 1029.1609, 1029.1268, 1029.079, 1029.0278, 1028.9784, 1028.9316, 1028.8855, 1028.8438, 1028.7987, 1028.7512, 1028.7098, 1028.6681, 1028.6208, 1028.5736, 1028.5209, 1028.4769, 1028.4277, 1028.3812, 1028.3267, 1028.2778, 1028.2312, 1028.1793, 1028.1226, 1028.0684, 1028.0138, 1027.9556, 1027.9081, 1027.8501, 1027.805, 1027.7501, 1027.6965, 1027.6437, 1027.5859, 1027.538, 1027.4825, 1027.4305, 1027.3748, 1027.3154, 1027.2516, 1027.1827, 1027.1165, 1027.0573, 1027.004, 1026.9536, 1026.8947, 1026.8308, 1026.757, 1026.6835, 1026.5898, 1026.4901, 1026.3896, 1026.2728, 1026.1797, 1026.0436, 1025.8846, 1025.7325, 1025.5847, 1025.4337, 1025.3278, 1025.209, 1025.1234, 1025.0189, 1024.8965, 1024.8118, 1024.495, 1024.112, 1023.98096, 1023.90704, 1023.8651, 1023.8391, 1023.82434, NaN, NaN, 1029.1846, 1029.1606, 1029.1226, 1029.0762, 1029.0269, 1028.9769, 1028.9347, 1028.886, 1028.837, 1028.789, 1028.7444, 1028.6996, 1028.647, 1028.6002, 1028.5535, 1028.4989, 1028.4458, 1028.3945, 1028.34, 1028.2812, 1028.229, 1028.1763, 1028.1265, 1028.0768, 1028.023, 1027.9711, 1027.9125, 1027.8604, 1027.8077, 1027.7504, 1027.7014, 1027.6444, 1027.5975, 1027.5356, 1027.4808, 1027.4263, 1027.3698, 1027.3021, 1027.2372, 1027.183, 1027.1333, 1027.071, 1026.9944, 1026.9382, 1026.8722, 1026.7993, 1026.7301, 1026.6495, 1026.5502, 1026.4524, 1026.3785, 1026.2886, 1026.1884, 1026.0646, 1025.9614, 1025.7906, 1025.6406, 1025.5121, 1025.3969, 1025.2496, 1025.0679, 1024.9209, 1024.6776, 1024.3029, 1024.1411, 1024.0469, 1023.9209, 1023.8457, 1023.8201, 1023.8026, NaN, NaN, 1029.2035, 1029.1758, 1029.139, 1029.0895, 1029.0433, 1028.9908, 1028.9463, 1028.893, 1028.8469, 1028.7971, 1028.7532, 1028.7069, 1028.6593, 1028.6129, 1028.567, 1028.5205, 1028.4783, 1028.4332, 1028.3867, 1028.3395, 1028.2976, 1028.2479, 1028.1947, 1028.1475, 1028.0996, 1028.0504, 1027.9965, 1027.9463, 1027.8926, 1027.8483, 1027.7986, 1027.7435, 1027.6912, 1027.6382, 1027.584, 1027.5355, 1027.4828, 1027.4143, 1027.357, 1027.3071, 1027.2556, 1027.1923, 1027.1405, 1027.091, 1027.03, 1026.9827, 1026.9327, 1026.8774, 1026.8206, 1026.727, 1026.6373, 1026.5618, 1026.4967, 1026.415, 1026.283, 1026.1768, 1026.0497, 1025.9028, 1025.773, 1025.6193, 1025.4492, 1025.302, 1025.1184, 1024.9758, 1024.816, 1024.3971, 1024.2657, 1024.1482, 1023.9527, 1023.849, 1023.82654, 1023.8104, NaN, NaN, 1029.2115, 1029.1843, 1029.1482, 1029.0988, 1029.0483, 1028.9995, 1028.9528, 1028.9059, 1028.8593, 1028.8088, 1028.7589, 1028.7091, 1028.669, 1028.6194, 1028.5675, 1028.5168, 1028.4656, 1028.4233, 1028.3752, 1028.3195, 1028.2637, 1028.201, 1028.1501, 1028.0942, 1028.0442, 1027.9945, 1027.9451, 1027.8925, 1027.8389, 1027.7789, 1027.7169, 1027.6584, 1027.5919, 1027.5386, 1027.4778, 1027.4109, 1027.3486, 1027.291, 1027.2294, 1027.17, 1027.0935, 1027.0128, 1026.9313, 1026.8567, 1026.7839, 1026.6815, 1026.5692, 1026.4823, 1026.3804, 1026.2114, 1026.1201, 1025.984, 1025.8447, 1025.6952, 1025.5568, 1025.4001, 1025.287, 1025.174, 1025.0332, 1024.9225, 1024.7639, 1024.4329, 1024.3055, 1024.2667, 1024.1091, 1023.85486, 1023.8289, 1023.8106, 1023.7985, NaN, NaN, 1029.1992, 1029.1719, 1029.1362, 1029.0852, 1029.0359, 1028.9913, 1028.9387, 1028.8857, 1028.8369, 1028.7828, 1028.7334, 1028.6887, 1028.6434, 1028.5957, 1028.5424, 1028.5027, 1028.4597, 1028.4144, 1028.3684, 1028.3221, 1028.2725, 1028.2292, 1028.1849, 1028.1438, 1028.0956, 1028.0516, 1028.0095, 1027.9618, 1027.912, 1027.864, 1027.8181, 1027.7759, 1027.7284, 1027.6874, 1027.6445, 1027.5988, 1027.5537, 1027.5143, 1027.472, 1027.4231, 1027.3651, 1027.3107, 1027.2622, 1027.2155, 1027.1605, 1027.1035, 1027.0338, 1026.9788, 1026.9186, 1026.8458, 1026.775, 1026.6971, 1026.5986, 1026.5078, 1026.3939, 1026.2756, 1026.12, 1025.9583, 1025.8202, 1025.6857, 1025.4929, 1025.3658, 1025.2295, 1025.124, 1025.017, 1024.8605, 1024.596, 1024.3927, 1024.3384, 1024.2064, 1023.9105, 1023.8728, 1023.84735, 1023.83344, NaN, NaN, 1029.2131, 1029.1882, 1029.1569, 1029.108, 1029.0591, 1029.0051, 1028.9531, 1028.9017, 1028.8539, 1028.8057, 1028.7493, 1028.697, 1028.6544, 1028.6117, 1028.563, 1028.5182, 1028.4697, 1028.4188, 1028.3672, 1028.3134, 1028.2655, 1028.2169, 1028.1678, 1028.1222, 1028.0797, 1028.0234, 1027.9736, 1027.9231, 1027.8789, 1027.829, 1027.7687, 1027.7079, 1027.6511, 1027.6013, 1027.5464, 1027.5005, 1027.4502, 1027.3997, 1027.342, 1027.2802, 1027.2147, 1027.1432, 1027.0688, 1027.0093, 1026.944, 1026.878, 1026.8279, 1026.7598, 1026.6787, 1026.5858, 1026.4728, 1026.3917, 1026.306, 1026.1726, 1026.0299, 1025.9031, 1025.7429, 1025.5896, 1025.4093, 1025.2844, 1025.1753, 1025.0487, 1024.9415, 1024.783, 1024.4735, 1024.2312, 1024.0505, 1023.91534, 1023.8981, NaN, NaN, 1029.2388, 1029.2098, 1029.1746, 1029.1261, 1029.074, 1029.0234, 1028.9716, 1028.9249, 1028.8745, 1028.8201, 1028.7625, 1028.7106, 1028.6577, 1028.6042, 1028.5587, 1028.5063, 1028.4595, 1028.4133, 1028.3627, 1028.3159, 1028.2672, 1028.2242, 1028.1722, 1028.1184, 1028.0706, 1028.0193, 1027.9668, 1027.9125, 1027.8575, 1027.8082, 1027.7571, 1027.7017, 1027.644, 1027.588, 1027.5398, 1027.4852, 1027.4409, 1027.3903, 1027.3315, 1027.2695, 1027.207, 1027.1445, 1027.07, 1027.0223, 1026.9651, 1026.8947, 1026.8118, 1026.7528, 1026.6677, 1026.5729, 1026.4978, 1026.3877, 1026.2588, 1026.137, 1025.9847, 1025.8384, 1025.6975, 1025.5507, 1025.354, 1025.2184, 1025.1166, 1024.9905, 1024.8035, 1024.4907, 1024.3416, 1024.2168, 1024.1437, 1024.0427, 1023.98535, 1023.9538, 1023.9349, NaN, NaN, 1029.2324, 1029.2007, 1029.1624, 1029.1077, 1029.0514, 1028.9966, 1028.9415, 1028.8912, 1028.8418, 1028.7844, 1028.7327, 1028.685, 1028.6322, 1028.5835, 1028.5316, 1028.4805, 1028.4296, 1028.3804, 1028.3331, 1028.2838, 1028.2312, 1028.183, 1028.1296, 1028.0773, 1028.025, 1027.9788, 1027.9247, 1027.868, 1027.813, 1027.7665, 1027.7151, 1027.6561, 1027.6069, 1027.5479, 1027.4893, 1027.4276, 1027.3691, 1027.3088, 1027.2533, 1027.1954, 1027.1201, 1027.0525, 1026.9756, 1026.8965, 1026.8271, 1026.748, 1026.6649, 1026.5742, 1026.4648, 1026.3185, 1026.1881, 1026.0813, 1025.9507, 1025.8254, 1025.65, 1025.496, 1025.3462, 1025.2196, 1025.0212, 1024.706, 1024.4468, 1024.2462, 1024.0782, 1024.0236, 1023.9396, 1023.81305, 1023.7582, 1023.73566, NaN, NaN, 1029.2223, 1029.1932, 1029.1547, 1029.1029, 1029.0532, 1029.0039, 1028.9526, 1028.9004, 1028.8506, 1028.798, 1028.7452, 1028.6914, 1028.6356, 1028.5863, 1028.5343, 1028.4836, 1028.4305, 1028.3826, 1028.3363, 1028.2865, 1028.2283, 1028.1769, 1028.1302, 1028.0785, 1028.0231, 1027.9651, 1027.9088, 1027.8694, 1027.8243, 1027.777, 1027.7289, 1027.6798, 1027.6246, 1027.568, 1027.5103, 1027.4552, 1027.4067, 1027.3542, 1027.3024, 1027.252, 1027.198, 1027.1467, 1027.0742, 1027.0192, 1026.9342, 1026.8597, 1026.7986, 1026.7163, 1026.6113, 1026.5203, 1026.4026, 1026.283, 1026.184, 1026.0575, 1025.897, 1025.7615, 1025.6702, 1025.501, 1025.3323, 1025.2222, 1025.0558, 1024.746, 1024.5057, 1024.1586, 1023.9754, 1023.80817, 1023.7262, 1023.6932, 1023.67694, NaN, NaN, 1029.2427, 1029.2188, 1029.184, 1029.13, 1029.0773, 1029.0216, 1028.9735, 1028.9252, 1028.8795, 1028.8331, 1028.7854, 1028.7388, 1028.6876, 1028.6388, 1028.5884, 1028.5392, 1028.4905, 1028.4453, 1028.4017, 1028.3574, 1028.308, 1028.2598, 1028.2073, 1028.1538, 1028.104, 1028.056, 1028.0099, 1027.9624, 1027.9053, 1027.8542, 1027.8048, 1027.7616, 1027.7133, 1027.6506, 1027.5956, 1027.5483, 1027.4987, 1027.4432, 1027.386, 1027.3363, 1027.2832, 1027.2252, 1027.1667, 1027.095, 1027.0331, 1026.9717, 1026.9227, 1026.8676, 1026.7898, 1026.696, 1026.5934, 1026.4956, 1026.4054, 1026.2456, 1026.1011, 1025.9668, 1025.8379, 1025.7377, 1025.556, 1025.3822, 1025.1526, 1024.936, 1024.6232, 1024.0249, 1023.7941, 1023.7431, 1023.7208, 1023.7018, 1023.6867, 1023.66406, 1023.65106, NaN, NaN, 1029.2301, 1029.2032, 1029.1683, 1029.1287, 1029.0874, 1029.047, 1028.9999, 1028.9548, 1028.9154, 1028.8724, 1028.8275, 1028.7837, 1028.7429, 1028.6951, 1028.6527, 1028.6097, 1028.5726, 1028.5325, 1028.4866, 1028.4436, 1028.4001, 1028.3545, 1028.3083, 1028.2659, 1028.2191, 1028.1771, 1028.133, 1028.0917, 1028.0499, 1028.0007, 1027.9562, 1027.908, 1027.863, 1027.8164, 1027.7736, 1027.7281, 1027.679, 1027.6349, 1027.5917, 1027.5471, 1027.5029, 1027.4525, 1027.403, 1027.3501, 1027.3008, 1027.2362, 1027.1711, 1027.1119, 1027.0499, 1026.989, 1026.9216, 1026.8473, 1026.7922, 1026.7274, 1026.6499, 1026.5645, 1026.4865, 1026.4059, 1026.2966, 1026.1774, 1026.084, 1025.9952, 1025.8945, 1025.7615, 1025.6602, 1025.5579, 1025.434, 1025.2721, 1025.0321, 1024.6802, 1024.1909, 1023.90576, 1023.71893, 1023.7022, 1023.6812, 1023.6644, 1023.6408, 1023.6345, NaN, NaN, 1029.2263, 1029.196, 1029.1602, 1029.1136, 1029.0632, 1029.0115, 1028.9581, 1028.9037, 1028.8512, 1028.8015, 1028.7432, 1028.6906, 1028.6421, 1028.5922, 1028.5438, 1028.4868, 1028.4397, 1028.3912, 1028.3384, 1028.2852, 1028.2295, 1028.17, 1028.118, 1028.0665, 1028.0269, 1027.9758, 1027.929, 1027.8785, 1027.8313, 1027.7778, 1027.7289, 1027.6797, 1027.6262, 1027.5759, 1027.5104, 1027.4583, 1027.4102, 1027.3491, 1027.2786, 1027.2134, 1027.1512, 1027.0919, 1027.0404, 1026.9851, 1026.8955, 1026.8197, 1026.7478, 1026.6526, 1026.5243, 1026.4248, 1026.2747, 1026.1482, 1026.0503, 1025.9146, 1025.785, 1025.6584, 1025.4681, 1025.3264, 1025.1619, 1024.8667, 1024.0447, 1023.75684, 1023.6872, 1023.6669, 1023.6494, 1023.63434, 1023.62164, NaN, NaN, 1029.2301, 1029.2036, 1029.1672, 1029.1155, 1029.0687, 1029.0234, 1028.9781, 1028.9304, 1028.8864, 1028.8291, 1028.7843, 1028.7318, 1028.6815, 1028.63, 1028.5815, 1028.5317, 1028.4805, 1028.4329, 1028.3805, 1028.328, 1028.2772, 1028.2286, 1028.178, 1028.1244, 1028.0712, 1028.0238, 1027.9745, 1027.9349, 1027.8859, 1027.8367, 1027.7795, 1027.722, 1027.6674, 1027.6176, 1027.5632, 1027.5137, 1027.4689, 1027.4185, 1027.3601, 1027.2976, 1027.2388, 1027.1941, 1027.1482, 1027.0944, 1027.0431, 1026.9712, 1026.8921, 1026.8259, 1026.7539, 1026.6521, 1026.5511, 1026.4435, 1026.3514, 1026.2683, 1026.1648, 1026.0779, 1025.9557, 1025.8591, 1025.7251, 1025.6184, 1025.4772, 1025.2968, 1024.9604, 1023.9557, 1023.8383, 1023.8185, 1023.7886, 1023.7575, 1023.713, 1023.6976, 1023.68463, NaN, NaN, 1029.2344, 1029.2079, 1029.1676, 1029.1128, 1029.0598, 1029.0078, 1028.9569, 1028.9069, 1028.8564, 1028.806, 1028.7513, 1028.7053, 1028.6592, 1028.6144, 1028.567, 1028.5216, 1028.4725, 1028.4231, 1028.3711, 1028.3229, 1028.2734, 1028.2214, 1028.17, 1028.1184, 1028.0682, 1028.0205, 1027.9537, 1027.8966, 1027.8436, 1027.7954, 1027.7324, 1027.6862, 1027.6426, 1027.5883, 1027.5284, 1027.4768, 1027.4207, 1027.3748, 1027.3242, 1027.2712, 1027.2177, 1027.1569, 1027.1, 1027.0254, 1026.9551, 1026.8921, 1026.8064, 1026.7166, 1026.5967, 1026.4846, 1026.3517, 1026.2294, 1026.1184, 1026.011, 1025.9103, 1025.7959, 1025.6582, 1025.4818, 1025.23, 1024.914, 1024.357, 1023.87463, 1023.85175, 1023.82996, 1023.808, 1023.7825, 1023.7581, 1023.73566, NaN, NaN, 1029.2421, 1029.2152, 1029.1782, 1029.1259, 1029.0781, 1029.0267, 1028.9751, 1028.9259, 1028.8733, 1028.8185, 1028.7683, 1028.7177, 1028.669, 1028.6189, 1028.5712, 1028.5223, 1028.4614, 1028.4081, 1028.3517, 1028.3038, 1028.2566, 1028.2062, 1028.1599, 1028.1149, 1028.0704, 1028.0304, 1027.9731, 1027.92, 1027.8729, 1027.8282, 1027.7766, 1027.7306, 1027.6798, 1027.6262, 1027.5731, 1027.5249, 1027.4742, 1027.434, 1027.3846, 1027.339, 1027.2749, 1027.2163, 1027.1644, 1027.1127, 1027.0444, 1026.9768, 1026.9154, 1026.8397, 1026.7568, 1026.6727, 1026.5874, 1026.4823, 1026.3712, 1026.2787, 1026.187, 1026.0736, 1025.9407, 1025.801, 1025.6493, 1025.5087, 1025.4, 1025.2555, 1024.9868, 1024.2039, 1023.8542, 1023.8398, 1023.82117, 1023.8007, 1023.77386, 1023.74835, 1023.7292, NaN, NaN, 1029.2463, 1029.2174, 1029.1802, 1029.1338, 1029.0972, 1029.0571, 1029.0154, 1028.9689, 1028.9225, 1028.8746, 1028.8314, 1028.7898, 1028.7433, 1028.701, 1028.6598, 1028.6196, 1028.577, 1028.5275, 1028.489, 1028.447, 1028.4, 1028.3527, 1028.3077, 1028.2646, 1028.2247, 1028.1777, 1028.1323, 1028.0857, 1028.0421, 1027.9867, 1027.9396, 1027.8861, 1027.8324, 1027.7827, 1027.7416, 1027.6981, 1027.6583, 1027.6068, 1027.5624, 1027.5168, 1027.4752, 1027.4307, 1027.3826, 1027.3286, 1027.2754, 1027.2114, 1027.1536, 1027.0775, 1027.0114, 1026.9454, 1026.8772, 1026.8008, 1026.7291, 1026.6519, 1026.5262, 1026.4269, 1026.342, 1026.2417, 1026.1748, 1026.0634, 1025.9681, 1025.8429, 1025.7148, 1025.5903, 1025.4862, 1025.3141, 1025.0715, 1024.6117, 1024.0472, 1023.8556, 1023.76276, 1023.6787, 1023.6567, 1023.63043, 1023.60736, 1023.57416, NaN, NaN, 1029.2473, 1029.2178, 1029.1765, 1029.1205, 1029.0725, 1029.0187, 1028.967, 1028.9142, 1028.8641, 1028.8124, 1028.7612, 1028.7114, 1028.6648, 1028.6138, 1028.5657, 1028.5121, 1028.4578, 1028.4025, 1028.3483, 1028.2865, 1028.2339, 1028.1809, 1028.1287, 1028.0807, 1028.0266, 1027.9706, 1027.9185, 1027.8667, 1027.8113, 1027.7488, 1027.6964, 1027.6367, 1027.5881, 1027.532, 1027.4757, 1027.4198, 1027.3715, 1027.2999, 1027.247, 1027.1917, 1027.1279, 1027.07, 1026.9897, 1026.9269, 1026.8606, 1026.7628, 1026.6671, 1026.5754, 1026.4651, 1026.3499, 1026.2576, 1026.1243, 1025.9878, 1025.895, 1025.8226, 1025.7104, 1025.5859, 1025.4183, 1025.1667, 1024.8901, 1024.5973, 1024.2378, 1023.8645, 1023.7269, 1023.64703, 1023.6064, 1023.56165, 1023.5111, NaN, NaN, 1029.2323, 1029.2035, 1029.1691, 1029.1191, 1029.0706, 1029.0199, 1028.9688, 1028.9125, 1028.8586, 1028.8025, 1028.7461, 1028.6902, 1028.639, 1028.5879, 1028.536, 1028.4885, 1028.4337, 1028.3787, 1028.3235, 1028.271, 1028.213, 1028.1632, 1028.1067, 1028.0483, 1027.9945, 1027.9382, 1027.8767, 1027.8228, 1027.7727, 1027.7227, 1027.669, 1027.6116, 1027.5548, 1027.5032, 1027.4478, 1027.3888, 1027.3348, 1027.2711, 1027.2188, 1027.1481, 1027.0845, 1027.0148, 1026.9336, 1026.8527, 1026.7897, 1026.7106, 1026.6133, 1026.5067, 1026.3699, 1026.285, 1026.1671, 1026.0353, 1025.9012, 1025.7513, 1025.6298, 1025.4734, 1025.3517, 1025.1589, 1024.7839, 1024.2107, 1023.80615, 1023.7799, 1023.7267, 1023.637, 1023.566, 1023.50903, NaN, NaN, 1029.2252, 1029.1967, 1029.161, 1029.1077, 1029.0537, 1029.0055, 1028.9572, 1028.903, 1028.8522, 1028.804, 1028.7546, 1028.7073, 1028.6589, 1028.6117, 1028.559, 1028.5131, 1028.4683, 1028.4264, 1028.3772, 1028.3287, 1028.2872, 1028.2362, 1028.1831, 1028.1266, 1028.0708, 1028.0195, 1027.9635, 1027.9102, 1027.8572, 1027.8068, 1027.7568, 1027.7034, 1027.6497, 1027.5986, 1027.5472, 1027.4967, 1027.4436, 1027.3909, 1027.343, 1027.2773, 1027.216, 1027.166, 1027.1134, 1027.0535, 1026.9922, 1026.9141, 1026.8241, 1026.7264, 1026.6577, 1026.5923, 1026.5135, 1026.4149, 1026.3107, 1026.184, 1026.0848, 1025.9565, 1025.8883, 1025.7498, 1025.6202, 1025.4949, 1025.3158, 1025.2147, 1025.0874, 1024.7502, 1024.1405, 1023.83203, 1023.79694, 1023.7536, 1023.69434, 1023.6507, 1023.62366, NaN, NaN, 1029.2262, 1029.2008, 1029.1664, 1029.1146, 1029.0638, 1029.0117, 1028.9589, 1028.9121, 1028.8625, 1028.8152, 1028.7595, 1028.7075, 1028.658, 1028.607, 1028.5585, 1028.5126, 1028.4681, 1028.4185, 1028.3671, 1028.3221, 1028.2819, 1028.2339, 1028.1892, 1028.1346, 1028.0846, 1028.0375, 1027.9888, 1027.9403, 1027.8893, 1027.849, 1027.7969, 1027.7427, 1027.6716, 1027.6128, 1027.5598, 1027.5101, 1027.449, 1027.3942, 1027.3524, 1027.3031, 1027.2454, 1027.1836, 1027.1144, 1027.0408, 1026.9795, 1026.9097, 1026.8296, 1026.7377, 1026.6412, 1026.5509, 1026.4417, 1026.3414, 1026.2405, 1026.1646, 1026.0426, 1025.9365, 1025.7449, 1025.6146, 1025.5018, 1025.3568, 1025.1744, 1025.0278, 1024.818, 1024.5515, 1024.3231, 1024.2239, 1024.0079, 1023.8473, 1023.69574, 1023.647, 1023.62274, 1023.6068, NaN, NaN, 1029.2198, 1029.1953, 1029.1602, 1029.1106, 1029.0624, 1029.013, 1028.9664, 1028.9198, 1028.8688, 1028.8179, 1028.768, 1028.7223, 1028.68, 1028.6278, 1028.5835, 1028.5327, 1028.4836, 1028.4313, 1028.3737, 1028.3202, 1028.2773, 1028.2288, 1028.1823, 1028.1327, 1028.0836, 1028.0397, 1027.9824, 1027.9335, 1027.8763, 1027.8259, 1027.7716, 1027.7198, 1027.6615, 1027.6044, 1027.5459, 1027.4872, 1027.4275, 1027.3682, 1027.3187, 1027.2604, 1027.2148, 1027.1592, 1027.0825, 1027.0138, 1026.9468, 1026.8807, 1026.8038, 1026.7222, 1026.6509, 1026.5951, 1026.5002, 1026.4004, 1026.2678, 1026.1111, 1025.9806, 1025.8561, 1025.6694, 1025.485, 1025.3441, 1025.1923, 1025.025, 1024.8091, 1024.6016, 1024.3674, 1024.2825, 1024.1536, 1023.91547, 1023.7846, 1023.6981, 1023.6776, NaN, NaN, 1029.2097, 1029.1809, 1029.1451, 1029.0969, 1029.055, 1029.0105, 1028.9619, 1028.9152, 1028.8694, 1028.8268, 1028.7843, 1028.7438, 1028.6946, 1028.6494, 1028.6036, 1028.557, 1028.5098, 1028.4615, 1028.4155, 1028.3756, 1028.3276, 1028.2891, 1028.2361, 1028.1748, 1028.1205, 1028.07, 1028.0157, 1027.9675, 1027.9167, 1027.8705, 1027.8282, 1027.7822, 1027.7325, 1027.6843, 1027.6356, 1027.583, 1027.5275, 1027.4683, 1027.4193, 1027.3717, 1027.3231, 1027.267, 1027.209, 1027.1322, 1027.0801, 1027.017, 1026.954, 1026.8987, 1026.8418, 1026.7682, 1026.6993, 1026.605, 1026.5134, 1026.4103, 1026.3097, 1026.2334, 1026.0808, 1025.9675, 1025.8372, 1025.7203, 1025.5674, 1025.416, 1025.263, 1025.1263, 1024.9991, 1024.8341, 1024.669, 1024.4117, 1024.3289, 1024.2717, 1024.2059, 1023.99457, 1023.82654, 1023.8024, NaN, NaN, 1029.182, 1029.1531, 1029.1211, 1029.0645, 1029.0117, 1028.9617, 1028.9094, 1028.858, 1028.7993, 1028.7444, 1028.6898, 1028.6343, 1028.5786, 1028.5227, 1028.4672, 1028.41, 1028.3423, 1028.2843, 1028.2334, 1028.1763, 1028.124, 1028.0667, 1028.0137, 1027.9541, 1027.9016, 1027.8502, 1027.7959, 1027.7319, 1027.6771, 1027.6191, 1027.5608, 1027.5066, 1027.4437, 1027.3688, 1027.3096, 1027.2548, 1027.191, 1027.1227, 1027.0663, 1027.004, 1026.9381, 1026.8687, 1026.8224, 1026.7552, 1026.6992, 1026.6389, 1026.557, 1026.4578, 1026.3414, 1026.2079, 1026.065, 1025.9218, 1025.7174, 1025.5424, 1025.3975, 1025.2546, 1025.1393, 1025.0056, 1024.8091, 1024.4932, 1024.3687, 1024.3131, 1024.2498, 1024.1722, 1024.0521, 1023.95856, NaN, NaN, 1029.2004, 1029.1754, 1029.145, 1029.1034, 1029.0609, 1029.0175, 1028.9679, 1028.9202, 1028.8806, 1028.8298, 1028.7793, 1028.735, 1028.6835, 1028.6362, 1028.5817, 1028.5377, 1028.4906, 1028.4359, 1028.3835, 1028.3337, 1028.2743, 1028.2174, 1028.1669, 1028.1221, 1028.0769, 1028.0215, 1027.9637, 1027.9124, 1027.8638, 1027.8118, 1027.7515, 1027.6924, 1027.6353, 1027.5785, 1027.5267, 1027.479, 1027.4233, 1027.3641, 1027.3135, 1027.2507, 1027.1774, 1027.119, 1027.0543, 1026.9968, 1026.9259, 1026.8657, 1026.7974, 1026.7174, 1026.6332, 1026.5529, 1026.4847, 1026.3964, 1026.2789, 1026.1567, 1026.0244, 1025.8391, 1025.6422, 1025.4628, 1025.3617, 1025.2473, 1025.0927, 1024.938, 1024.7792, 1024.4255, 1024.2983, 1024.2361, 1024.1575, 1023.9747, 1023.8047, 1023.71124, NaN, NaN, 1029.192, 1029.1669, 1029.1385, 1029.0989, 1029.0597, 1029.0148, 1028.9648, 1028.9246, 1028.8801, 1028.8376, 1028.7935, 1028.7479, 1028.7065, 1028.659, 1028.6116, 1028.5632, 1028.5189, 1028.4741, 1028.4294, 1028.3811, 1028.3379, 1028.2914, 1028.2384, 1028.1929, 1028.1495, 1028.1033, 1028.0496, 1028.0016, 1027.9567, 1027.9064, 1027.8656, 1027.8209, 1027.7771, 1027.7295, 1027.6868, 1027.6481, 1027.5947, 1027.546, 1027.4938, 1027.4507, 1027.402, 1027.3448, 1027.291, 1027.2369, 1027.1864, 1027.1406, 1027.0992, 1027.0514, 1027.0029, 1026.9503, 1026.8969, 1026.853, 1026.7998, 1026.7516, 1026.7031, 1026.6454, 1026.5856, 1026.4917, 1026.3906, 1026.3147, 1026.235, 1026.1338, 1026.0632, 1025.9794, 1025.7787, 1025.6365, 1025.5696, 1025.462, 1025.3284, 1025.1774, 1025.049, 1024.8909, 1024.7482, 1024.4167, 1024.2562, 1024.0128, 1023.9509, 1023.8147, 1023.74, 1023.69745, NaN, NaN, 1029.1744, 1029.1497, 1029.1134, 1029.0653, 1029.0181, 1028.9741, 1028.929, 1028.8896, 1028.8469, 1028.8036, 1028.755, 1028.7067, 1028.652, 1028.6058, 1028.5518, 1028.4893, 1028.4294, 1028.3708, 1028.3048, 1028.2389, 1028.1826, 1028.1279, 1028.06, 1028.0054, 1027.939, 1027.8777, 1027.8162, 1027.765, 1027.7158, 1027.6595, 1027.6018, 1027.5283, 1027.4543, 1027.3885, 1027.3339, 1027.2793, 1027.2216, 1027.1696, 1027.1119, 1027.0535, 1026.9994, 1026.936, 1026.8837, 1026.8326, 1026.7854, 1026.7201, 1026.6482, 1026.562, 1026.4834, 1026.3861, 1026.2898, 1026.1913, 1026.0277, 1025.8518, 1025.6971, 1025.5117, 1025.3671, 1025.2451, 1025.1089, 1024.9603, 1024.741, 1024.3416, 1024.0161, 1023.8838, 1023.79346, 1023.7566, 1023.6856, NaN, NaN, 1029.1692, 1029.1427, 1029.1067, 1029.0624, 1029.0193, 1028.9786, 1028.9355, 1028.8921, 1028.8486, 1028.8048, 1028.7606, 1028.7152, 1028.666, 1028.6201, 1028.5745, 1028.5269, 1028.4758, 1028.4233, 1028.3743, 1028.3181, 1028.2625, 1028.201, 1028.1417, 1028.0828, 1028.0325, 1027.9742, 1027.925, 1027.8684, 1027.8033, 1027.7375, 1027.6691, 1027.6053, 1027.551, 1027.4867, 1027.4288, 1027.3672, 1027.3044, 1027.2437, 1027.1838, 1027.133, 1027.0844, 1027.0392, 1026.9934, 1026.9341, 1026.8678, 1026.8097, 1026.7512, 1026.6829, 1026.6034, 1026.499, 1026.4147, 1026.3171, 1026.1815, 1026.0497, 1025.908, 1025.7637, 1025.6163, 1025.4468, 1025.3005, 1025.21, 1025.0631, 1024.8735, 1024.6976, 1024.504, 1024.0001, 1023.8848, 1023.8632, 1023.8416, 1023.8107, 1023.7485, 1023.6697, NaN, NaN, 1029.1755, 1029.15, 1029.1144, 1029.0703, 1029.0214, 1028.973, 1028.923, 1028.8728, 1028.8184, 1028.7623, 1028.7045, 1028.6505, 1028.5973, 1028.5408, 1028.4891, 1028.4355, 1028.3871, 1028.337, 1028.2814, 1028.225, 1028.1692, 1028.1189, 1028.0659, 1028.0128, 1027.9519, 1027.89, 1027.8307, 1027.784, 1027.7233, 1027.647, 1027.5792, 1027.5167, 1027.4532, 1027.391, 1027.3378, 1027.2742, 1027.2101, 1027.1483, 1027.0984, 1027.0518, 1026.9996, 1026.9514, 1026.9044, 1026.8397, 1026.7753, 1026.702, 1026.6434, 1026.5668, 1026.4697, 1026.3052, 1026.1919, 1026.0151, 1025.7798, 1025.6061, 1025.4385, 1025.3528, 1025.2024, 1025.0825, 1024.9856, 1024.8121, 1024.252, 1023.89185, 1023.86487, 1023.83154, 1023.7938, 1023.7157, 1023.6681, NaN, NaN, 1029.1859, 1029.1592, 1029.1224, 1029.0802, 1029.0339, 1028.9915, 1028.949, 1028.9058, 1028.8591, 1028.8123, 1028.7609, 1028.7092, 1028.6583, 1028.6123, 1028.5659, 1028.5173, 1028.4664, 1028.4185, 1028.3583, 1028.3077, 1028.2651, 1028.2206, 1028.17, 1028.1119, 1028.0581, 1028.0109, 1027.9504, 1027.8881, 1027.8334, 1027.765, 1027.699, 1027.6313, 1027.5682, 1027.4991, 1027.4369, 1027.3773, 1027.3109, 1027.2369, 1027.1758, 1027.1171, 1027.0726, 1027.0251, 1026.975, 1026.916, 1026.8613, 1026.8015, 1026.7229, 1026.6752, 1026.636, 1026.5957, 1026.5002, 1026.3762, 1026.3038, 1026.1583, 1026.0826, 1025.9019, 1025.7396, 1025.5543, 1025.4001, 1025.2905, 1025.1554, 1024.9641, 1024.6863, 1023.94434, 1023.87823, 1023.795, 1023.7062, 1023.6709, 1023.6547, 1023.6381, NaN, NaN, 1029.163, 1029.1376, 1029.1025, 1029.051, 1029.0067, 1028.9601, 1028.9132, 1028.8599, 1028.8119, 1028.7528, 1028.6951, 1028.6426, 1028.5885, 1028.535, 1028.4845, 1028.43, 1028.3744, 1028.3175, 1028.267, 1028.2262, 1028.1759, 1028.1276, 1028.0834, 1028.0372, 1027.9893, 1027.929, 1027.8667, 1027.7933, 1027.7247, 1027.661, 1027.5695, 1027.4823, 1027.4067, 1027.3383, 1027.2671, 1027.2115, 1027.1583, 1027.1019, 1027.0377, 1026.9803, 1026.934, 1026.8827, 1026.8291, 1026.7761, 1026.7246, 1026.662, 1026.5891, 1026.5106, 1026.3997, 1026.3008, 1026.1891, 1026.0353, 1025.8595, 1025.6024, 1025.3729, 1025.2285, 1025.1212, 1025.0234, 1024.7526, 1024.269, 1023.81433, 1023.74274, 1023.71277, 1023.69086, 1023.67163, NaN, NaN, 1029.1683, 1029.1437, 1029.1108, 1029.0565, 1029.003, 1028.9496, 1028.8994, 1028.849, 1028.7982, 1028.7499, 1028.6964, 1028.6483, 1028.5973, 1028.5481, 1028.5051, 1028.4624, 1028.4188, 1028.3776, 1028.322, 1028.279, 1028.2318, 1028.1865, 1028.1423, 1028.0985, 1028.0514, 1028.0049, 1027.9569, 1027.8988, 1027.8243, 1027.744, 1027.6542, 1027.5494, 1027.4735, 1027.4015, 1027.3326, 1027.2783, 1027.2218, 1027.1649, 1027.1145, 1027.0677, 1027.0198, 1026.972, 1026.9165, 1026.8651, 1026.8134, 1026.7678, 1026.7201, 1026.6683, 1026.5908, 1026.5232, 1026.4346, 1026.3296, 1026.1858, 1026.0098, 1025.8589, 1025.7389, 1025.5248, 1025.2971, 1025.1311, 1024.8934, 1024.543, 1023.9742, 1023.85657, 1023.8282, 1023.73846, 1023.6863, 1023.65955, 1023.64105, NaN, NaN, 1029.1721, 1029.1488, 1029.114, 1029.0701, 1029.0253, 1028.977, 1028.9279, 1028.878, 1028.8307, 1028.7769, 1028.7256, 1028.677, 1028.6266, 1028.5831, 1028.536, 1028.4905, 1028.4456, 1028.4072, 1028.3666, 1028.3151, 1028.2695, 1028.226, 1028.1792, 1028.1417, 1028.0887, 1028.0375, 1027.9928, 1027.9406, 1027.8735, 1027.7782, 1027.667, 1027.5948, 1027.5266, 1027.4746, 1027.4222, 1027.3702, 1027.3029, 1027.2446, 1027.1945, 1027.15, 1027.1091, 1027.0659, 1027.0278, 1026.978, 1026.937, 1026.8953, 1026.8513, 1026.8102, 1026.7717, 1026.7278, 1026.6821, 1026.629, 1026.5845, 1026.5353, 1026.4379, 1026.2926, 1026.0813, 1025.912, 1025.6768, 1025.4646, 1025.2814, 1025.1235, 1024.9636, 1024.8044, 1024.519, 1024.12, 1023.86774, 1023.7276, 1023.60065, 1023.5649, 1023.54083, 1023.52203, NaN, NaN, 1029.1742, 1029.1505, 1029.1166, 1029.0676, 1029.0194, 1028.962, 1028.9154, 1028.871, 1028.8188, 1028.7745, 1028.7241, 1028.662, 1028.6089, 1028.5569, 1028.5087, 1028.4619, 1028.4156, 1028.3685, 1028.3201, 1028.2686, 1028.2264, 1028.1744, 1028.129, 1028.0747, 1028.0326, 1027.9917, 1027.9379, 1027.8829, 1027.8209, 1027.76, 1027.6779, 1027.5598, 1027.489, 1027.4337, 1027.3838, 1027.3414, 1027.269, 1027.2179, 1027.1671, 1027.1267, 1027.0851, 1027.0449, 1026.9929, 1026.9427, 1026.8966, 1026.8512, 1026.8053, 1026.7549, 1026.704, 1026.6519, 1026.6025, 1026.5474, 1026.4691, 1026.329, 1026.0933, 1025.8833, 1025.6525, 1025.4153, 1025.3103, 1025.1287, 1024.9828, 1024.8129, 1024.2734, 1023.83704, 1023.61743, 1023.5688, 1023.54614, 1023.5231, 1023.50714, NaN, NaN, 1029.1648, 1029.1348, 1029.0996, 1029.0538, 1029.0049, 1028.9613, 1028.9122, 1028.864, 1028.8148, 1028.7736, 1028.723, 1028.6732, 1028.6262, 1028.5723, 1028.525, 1028.4791, 1028.4307, 1028.384, 1028.3372, 1028.2931, 1028.2482, 1028.1901, 1028.148, 1028.1023, 1028.0541, 1028.003, 1027.9442, 1027.8807, 1027.814, 1027.7482, 1027.666, 1027.5975, 1027.5424, 1027.4861, 1027.4308, 1027.3789, 1027.3119, 1027.2556, 1027.2133, 1027.1674, 1027.1223, 1027.0774, 1027.028, 1026.9764, 1026.925, 1026.882, 1026.8364, 1026.7924, 1026.7496, 1026.701, 1026.6426, 1026.5897, 1026.5468, 1026.498, 1026.4164, 1026.2278, 1026.0156, 1025.8556, 1025.628, 1025.3663, 1025.1707, 1025.011, 1024.9296, 1024.6467, 1023.7673, 1023.5951, 1023.5674, 1023.54333, 1023.5276, NaN, NaN, 1029.146, 1029.1238, 1029.0875, 1029.0367, 1028.9856, 1028.9407, 1028.8993, 1028.8523, 1028.7997, 1028.7483, 1028.7006, 1028.6577, 1028.6112, 1028.5637, 1028.521, 1028.471, 1028.425, 1028.3773, 1028.3307, 1028.2863, 1028.243, 1028.1935, 1028.1478, 1028.0984, 1028.0482, 1027.9966, 1027.9401, 1027.8722, 1027.8071, 1027.7407, 1027.6652, 1027.5989, 1027.5339, 1027.4598, 1027.3969, 1027.3264, 1027.2645, 1027.2059, 1027.1509, 1027.104, 1027.057, 1027.0013, 1026.9565, 1026.917, 1026.8768, 1026.8422, 1026.8016, 1026.7587, 1026.7192, 1026.6721, 1026.605, 1026.5503, 1026.4908, 1026.3938, 1026.2357, 1026.053, 1025.8859, 1025.65, 1025.5145, 1025.3447, 1025.2389, 1025.1165, 1025.0729, 1024.8708, 1024.5765, 1024.281, 1023.96094, 1023.81287, 1023.6472, 1023.5995, 1023.5644, 1023.5474, NaN, NaN, 1029.1654, 1029.1412, 1029.1075, 1029.0558, 1029.0059, 1028.9562, 1028.908, 1028.8588, 1028.8114, 1028.7651, 1028.714, 1028.6647, 1028.6174, 1028.571, 1028.5256, 1028.4756, 1028.4263, 1028.3704, 1028.3151, 1028.2675, 1028.2129, 1028.1642, 1028.1136, 1028.0591, 1027.9991, 1027.9415, 1027.8746, 1027.8052, 1027.7184, 1027.6418, 1027.5693, 1027.4945, 1027.418, 1027.3344, 1027.2748, 1027.216, 1027.151, 1027.09, 1027.0358, 1026.9893, 1026.942, 1026.8947, 1026.8417, 1026.7924, 1026.739, 1026.6736, 1026.613, 1026.5469, 1026.4559, 1026.3419, 1026.1749, 1026.03, 1025.788, 1025.5862, 1025.4491, 1025.3019, 1025.1875, 1025.0931, 1024.924, 1024.6984, 1024.2584, 1023.9711, 1023.8839, 1023.746, 1023.6898, 1023.673, NaN, NaN, 1029.1487, 1029.1237, 1029.0916, 1029.0482, 1029.0065, 1028.9586, 1028.9078, 1028.8635, 1028.8131, 1028.7632, 1028.7177, 1028.6677, 1028.6174, 1028.5691, 1028.5211, 1028.476, 1028.4244, 1028.3649, 1028.316, 1028.2662, 1028.2103, 1028.1642, 1028.1113, 1028.0586, 1027.9922, 1027.932, 1027.8629, 1027.8007, 1027.7308, 1027.6606, 1027.5901, 1027.5309, 1027.4698, 1027.3993, 1027.3423, 1027.2777, 1027.2228, 1027.1724, 1027.1194, 1027.0667, 1027.0195, 1026.97, 1026.9215, 1026.8778, 1026.8204, 1026.7654, 1026.702, 1026.648, 1026.5826, 1026.5106, 1026.4059, 1026.2875, 1026.158, 1026.0055, 1025.8025, 1025.6444, 1025.5242, 1025.3441, 1025.1886, 1025.0754, 1024.9276, 1024.7799, 1024.5243, 1024.2762, 1024.0846, 1023.87024, 1023.8037, 1023.7901, NaN, NaN, 1029.1677, 1029.1434, 1029.1094, 1029.0646, 1029.0184, 1028.9723, 1028.9243, 1028.8759, 1028.8263, 1028.779, 1028.7303, 1028.6812, 1028.6338, 1028.5869, 1028.5371, 1028.4886, 1028.4376, 1028.3842, 1028.3301, 1028.2737, 1028.2211, 1028.1672, 1028.1158, 1028.0635, 1028.0054, 1027.945, 1027.8763, 1027.8087, 1027.7338, 1027.6709, 1027.5947, 1027.5294, 1027.4734, 1027.4104, 1027.3477, 1027.2937, 1027.2424, 1027.1902, 1027.1445, 1027.0999, 1027.0543, 1027.0094, 1026.9597, 1026.9102, 1026.8597, 1026.8097, 1026.7528, 1026.6895, 1026.626, 1026.5419, 1026.4299, 1026.3108, 1026.1776, 1026.0233, 1025.7766, 1025.6272, 1025.533, 1025.3938, 1025.2535, 1025.1377, 1025.0447, 1024.9355, 1024.744, 1024.3156, 1024.1367, 1024.0107, 1023.8475, 1023.80206, 1023.784, NaN, NaN, 1029.1576, 1029.1333, 1029.1023, 1029.0594, 1029.0208, 1028.9777, 1028.9354, 1028.8933, 1028.8527, 1028.8076, 1028.7603, 1028.7139, 1028.6683, 1028.6229, 1028.5775, 1028.5271, 1028.4778, 1028.4271, 1028.3739, 1028.3225, 1028.2661, 1028.2119, 1028.1595, 1028.108, 1028.0598, 1028.0023, 1027.9478, 1027.8921, 1027.8348, 1027.7657, 1027.7004, 1027.6505, 1027.6014, 1027.5435, 1027.4835, 1027.4241, 1027.3616, 1027.3156, 1027.2673, 1027.213, 1027.1635, 1027.1124, 1027.0652, 1027.0205, 1026.9783, 1026.9359, 1026.8853, 1026.8258, 1026.7687, 1026.706, 1026.6375, 1026.5531, 1026.4563, 1026.2983, 1026.1743, 1026.059, 1025.8602, 1025.6316, 1025.4669, 1025.2709, 1025.128, 1024.9955, 1024.8962, 1024.7458, 1024.4934, 1024.126, 1023.91504, 1023.81525, 1023.7751, NaN, NaN, 1029.145, 1029.1195, 1029.0857, 1029.0345, 1028.9829, 1028.9342, 1028.8871, 1028.8352, 1028.7844, 1028.7302, 1028.6758, 1028.623, 1028.5697, 1028.5166, 1028.4625, 1028.4126, 1028.3595, 1028.3021, 1028.2368, 1028.1843, 1028.1306, 1028.0801, 1028.0242, 1027.9714, 1027.9161, 1027.8605, 1027.8016, 1027.7487, 1027.6993, 1027.6406, 1027.5853, 1027.5325, 1027.4781, 1027.4261, 1027.3745, 1027.3235, 1027.2761, 1027.2295, 1027.1848, 1027.142, 1027.0912, 1027.0438, 1027.001, 1026.9556, 1026.9113, 1026.8514, 1026.7887, 1026.7283, 1026.6539, 1026.57, 1026.4425, 1026.3324, 1026.2253, 1026.0536, 1025.8256, 1025.6233, 1025.5044, 1025.3496, 1025.1732, 1025.0076, 1024.8411, 1024.6573, 1024.4689, 1024.2389, 1024.0206, 1023.9347, 1023.8607, 1023.8412, NaN, NaN, 1029.1492, 1029.1215, 1029.0884, 1029.0498, 1029.0139, 1028.9691, 1028.9237, 1028.8807, 1028.835, 1028.7948, 1028.755, 1028.712, 1028.6719, 1028.6276, 1028.5828, 1028.5383, 1028.4934, 1028.4467, 1028.4005, 1028.3567, 1028.308, 1028.2565, 1028.1981, 1028.1478, 1028.1024, 1028.0542, 1028.006, 1027.9518, 1027.9059, 1027.8431, 1027.7908, 1027.747, 1027.6931, 1027.6365, 1027.5867, 1027.5271, 1027.4681, 1027.4127, 1027.3625, 1027.3097, 1027.2576, 1027.2046, 1027.1523, 1027.1036, 1027.0526, 1027.0023, 1026.959, 1026.9082, 1026.8494, 1026.7993, 1026.7346, 1026.6631, 1026.5862, 1026.5011, 1026.4072, 1026.2792, 1026.1309, 1025.9117, 1025.7347, 1025.5848, 1025.4069, 1025.2306, 1025.124, 1025.0203, 1024.8887, 1024.7686, 1024.5468, 1024.1826, 1024.0707, 1023.9488, 1023.9311, NaN, NaN, 1029.1571, 1029.1313, 1029.0964, 1029.0533, 1029.0135, 1028.9673, 1028.9198, 1028.8761, 1028.832, 1028.7869, 1028.7405, 1028.6943, 1028.6447, 1028.6035, 1028.5591, 1028.5117, 1028.4639, 1028.4165, 1028.373, 1028.3282, 1028.2837, 1028.2301, 1028.1847, 1028.1362, 1028.0848, 1028.0294, 1027.9844, 1027.9243, 1027.8705, 1027.8135, 1027.76, 1027.6995, 1027.6418, 1027.5752, 1027.5234, 1027.4692, 1027.4022, 1027.3427, 1027.2941, 1027.2415, 1027.1915, 1027.1384, 1027.0939, 1027.0479, 1027.0007, 1026.9541, 1026.9015, 1026.8499, 1026.8031, 1026.7478, 1026.6853, 1026.6185, 1026.5297, 1026.4523, 1026.3247, 1026.167, 1026.0105, 1025.83, 1025.6753, 1025.5391, 1025.3936, 1025.2479, 1025.1235, 1025.0491, 1024.9805, 1024.847, 1024.7722, 1024.6646, 1024.5597, 1024.3468, 1023.939, 1023.78644, 1023.7678, 1023.7573, NaN, NaN, 1029.1614, 1029.135, 1029.1024, 1029.0491, 1028.9982, 1028.9484, 1028.8949, 1028.8455, 1028.7954, 1028.7422, 1028.6895, 1028.6354, 1028.5824, 1028.528, 1028.4634, 1028.4135, 1028.3545, 1028.298, 1028.2499, 1028.1941, 1028.1259, 1028.0717, 1028.0118, 1027.958, 1027.9019, 1027.8372, 1027.7782, 1027.7279, 1027.6727, 1027.6144, 1027.5461, 1027.4891, 1027.4243, 1027.3589, 1027.2935, 1027.2422, 1027.1833, 1027.1323, 1027.0769, 1027.0225, 1026.9767, 1026.9147, 1026.8618, 1026.814, 1026.7584, 1026.6906, 1026.597, 1026.4888, 1026.3759, 1026.265, 1026.129, 1025.9321, 1025.7273, 1025.5762, 1025.4703, 1025.3601, 1025.2689, 1025.0968, 1024.9313, 1024.7965, 1024.7043, 1024.6068, 1024.482, 1024.2108, 1023.9183, 1023.7907, 1023.7668, 1023.754, NaN, NaN, 1029.1713, 1029.147, 1029.1118, 1029.0625, 1029.0094, 1028.9603, 1028.9146, 1028.8674, 1028.8209, 1028.7697, 1028.7228, 1028.677, 1028.6288, 1028.5833, 1028.5267, 1028.4739, 1028.4172, 1028.3678, 1028.3137, 1028.2563, 1028.1962, 1028.1409, 1028.0807, 1028.0327, 1027.9756, 1027.916, 1027.8473, 1027.7753, 1027.7139, 1027.648, 1027.5851, 1027.5265, 1027.4767, 1027.4128, 1027.3552, 1027.305, 1027.2426, 1027.1869, 1027.1356, 1027.073, 1027.0172, 1026.959, 1026.8948, 1026.8282, 1026.7706, 1026.7084, 1026.6241, 1026.5254, 1026.4191, 1026.2972, 1026.1788, 1025.9957, 1025.7048, 1025.5209, 1025.3729, 1025.2651, 1025.0548, 1024.9423, 1024.8496, 1024.7288, 1024.6494, 1024.5686, 1024.3591, 1023.91486, 1023.7929, 1023.77, 1023.7468, NaN, NaN, 1029.1697, 1029.1454, 1029.1096, 1029.0603, 1029.0051, 1028.9531, 1028.905, 1028.856, 1028.8055, 1028.7571, 1028.7189, 1028.6675, 1028.616, 1028.564, 1028.5151, 1028.4567, 1028.4062, 1028.3563, 1028.304, 1028.249, 1028.196, 1028.1438, 1028.094, 1028.0448, 1027.9954, 1027.9386, 1027.8815, 1027.8319, 1027.7766, 1027.7173, 1027.6628, 1027.6069, 1027.5476, 1027.4888, 1027.4384, 1027.3906, 1027.334, 1027.2825, 1027.2281, 1027.1726, 1027.1234, 1027.0673, 1027.0106, 1026.9595, 1026.9054, 1026.8396, 1026.7694, 1026.7051, 1026.619, 1026.5236, 1026.4203, 1026.3141, 1026.2063, 1026.0543, 1025.8768, 1025.6666, 1025.4489, 1025.254, 1025.1088, 1024.951, 1024.8353, 1024.7734, 1024.687, 1024.6132, 1024.4962, 1023.932, 1023.79175, 1023.7573, 1023.732, NaN, NaN, 1029.1831, 1029.1561, 1029.1241, 1029.0797, 1029.0363, 1028.9889, 1028.9443, 1028.8949, 1028.8528, 1028.8044, 1028.7622, 1028.718, 1028.672, 1028.627, 1028.5809, 1028.5338, 1028.4866, 1028.4435, 1028.3958, 1028.3455, 1028.297, 1028.2471, 1028.2, 1028.1492, 1028.0977, 1028.0422, 1027.9929, 1027.9337, 1027.8881, 1027.838, 1027.7843, 1027.727, 1027.6832, 1027.6274, 1027.5667, 1027.5088, 1027.461, 1027.4053, 1027.3583, 1027.3016, 1027.2444, 1027.1921, 1027.1442, 1027.0979, 1027.0519, 1027.0077, 1026.9558, 1026.9021, 1026.8414, 1026.7856, 1026.7262, 1026.648, 1026.5708, 1026.465, 1026.3468, 1026.2434, 1026.1152, 1025.968, 1025.8467, 1025.6848, 1025.5466, 1025.3453, 1025.1854, 1025.0256, 1024.8217, 1024.7102, 1024.6442, 1024.5597, 1024.2833, 1023.9231, 1023.8376, 1023.7516, NaN, NaN, 1029.1763, 1029.1483, 1029.1118, 1029.061, 1029.0143, 1028.9644, 1028.9192, 1028.8701, 1028.82, 1028.7703, 1028.7213, 1028.674, 1028.6198, 1028.5724, 1028.5153, 1028.4598, 1028.4098, 1028.3596, 1028.3057, 1028.2474, 1028.188, 1028.1326, 1028.0762, 1028.0239, 1027.9667, 1027.9022, 1027.8359, 1027.7725, 1027.7152, 1027.652, 1027.5979, 1027.5345, 1027.4747, 1027.4159, 1027.3522, 1027.2826, 1027.2224, 1027.1661, 1027.0986, 1027.043, 1026.991, 1026.9401, 1026.8864, 1026.8257, 1026.7404, 1026.6538, 1026.5189, 1026.422, 1026.3168, 1026.1963, 1026.0472, 1025.8995, 1025.7365, 1025.5428, 1025.4354, 1025.2798, 1025.1069, 1024.9546, 1024.8342, 1024.7101, 1024.6062, 1024.3718, 1024.1425, 1024.0819, 1023.935, 1023.7736, 1023.75006, NaN, NaN, 1029.1794, 1029.1505, 1029.1177, 1029.0685, 1029.0231, 1028.9753, 1028.9269, 1028.8777, 1028.8314, 1028.7811, 1028.7352, 1028.6848, 1028.6368, 1028.5835, 1028.5269, 1028.4758, 1028.4305, 1028.3806, 1028.3301, 1028.2793, 1028.224, 1028.1677, 1028.1187, 1028.0638, 1028.0178, 1027.9642, 1027.9089, 1027.8516, 1027.7936, 1027.7311, 1027.6637, 1027.5996, 1027.5464, 1027.48, 1027.4172, 1027.3523, 1027.2905, 1027.235, 1027.174, 1027.1042, 1027.0413, 1026.9756, 1026.9144, 1026.8517, 1026.7819, 1026.7217, 1026.6476, 1026.5665, 1026.4463, 1026.2858, 1026.1469, 1025.9514, 1025.789, 1025.6614, 1025.5265, 1025.3491, 1025.1808, 1025.0754, 1025.0283, 1024.943, 1024.8013, 1024.6189, 1024.3984, 1024.1835, 1023.91547, 1023.8699, 1023.80664, 1023.7856, NaN, NaN, 1029.1896, 1029.1608, 1029.1215, 1029.0703, 1029.0181, 1028.9714, 1028.9177, 1028.8597, 1028.8134, 1028.7649, 1028.7109, 1028.6566, 1028.6062, 1028.5538, 1028.4993, 1028.4382, 1028.3795, 1028.3263, 1028.2668, 1028.206, 1028.1425, 1028.0911, 1028.032, 1027.9724, 1027.9215, 1027.8634, 1027.8081, 1027.7532, 1027.6991, 1027.6493, 1027.5859, 1027.5157, 1027.4583, 1027.3994, 1027.3402, 1027.2859, 1027.2235, 1027.1621, 1027.0916, 1027.0214, 1026.96, 1026.8967, 1026.8398, 1026.7751, 1026.7117, 1026.6469, 1026.5684, 1026.4885, 1026.3395, 1026.2008, 1026.0795, 1025.9396, 1025.8297, 1025.6188, 1025.3912, 1025.2867, 1025.1719, 1025.0354, 1024.9183, 1024.743, 1024.6052, 1024.4171, 1024.1296, 1023.9625, 1023.8959, 1023.85815, 1023.8325, NaN, NaN, 1029.1868, 1029.1573, 1029.1191, 1029.0673, 1029.0148, 1028.9662, 1028.9181, 1028.8702, 1028.8258, 1028.7709, 1028.7194, 1028.6669, 1028.6157, 1028.5686, 1028.5187, 1028.464, 1028.4082, 1028.3501, 1028.2916, 1028.2374, 1028.1774, 1028.1145, 1028.0629, 1028.0017, 1027.949, 1027.8955, 1027.8464, 1027.7914, 1027.7435, 1027.684, 1027.6309, 1027.5834, 1027.5309, 1027.4739, 1027.4047, 1027.3486, 1027.2817, 1027.2096, 1027.1366, 1027.0807, 1027.0215, 1026.9592, 1026.91, 1026.846, 1026.7761, 1026.707, 1026.6344, 1026.549, 1026.4702, 1026.3763, 1026.2361, 1026.068, 1025.9175, 1025.7474, 1025.6459, 1025.582, 1025.4459, 1025.3094, 1025.1434, 1025.0121, 1024.8901, 1024.7185, 1024.5698, 1024.4453, 1024.2147, 1023.9607, 1023.91345, 1023.8857, 1023.8691, 1023.85785, NaN, NaN, 1029.1975, 1029.1681, 1029.1279, 1029.0781, 1029.0214, 1028.9641, 1028.9106, 1028.8506, 1028.7933, 1028.7426, 1028.6963, 1028.6428, 1028.5966, 1028.5479, 1028.4976, 1028.4452, 1028.3904, 1028.3397, 1028.2864, 1028.2273, 1028.1759, 1028.1259, 1028.0714, 1028.0154, 1027.9613, 1027.8995, 1027.8439, 1027.7977, 1027.7428, 1027.6826, 1027.6237, 1027.5726, 1027.5187, 1027.4686, 1027.4185, 1027.3618, 1027.296, 1027.2314, 1027.1655, 1027.1138, 1027.0676, 1027.0013, 1026.9259, 1026.8491, 1026.777, 1026.7073, 1026.616, 1026.5508, 1026.4458, 1026.2981, 1026.1897, 1026.0323, 1025.882, 1025.7527, 1025.5916, 1025.3961, 1025.277, 1025.2002, 1025.1128, 1024.9832, 1024.8634, 1024.719, 1024.565, 1024.3972, 1024.0732, 1023.90753, 1023.8636, 1023.85504, NaN, NaN, 1029.1562, 1029.1302, 1029.092, 1029.0405, 1028.978, 1028.9205, 1028.863, 1028.8113, 1028.7606, 1028.7097, 1028.6593, 1028.607, 1028.5591, 1028.5066, 1028.4574, 1028.4082, 1028.3557, 1028.3035, 1028.2477, 1028.1958, 1028.141, 1028.0918, 1028.0381, 1027.9948, 1027.9481, 1027.8925, 1027.8348, 1027.7755, 1027.7155, 1027.6589, 1027.5941, 1027.5338, 1027.4674, 1027.4037, 1027.3438, 1027.2921, 1027.2316, 1027.1666, 1027.1033, 1027.0475, 1026.9763, 1026.9043, 1026.8237, 1026.7406, 1026.6462, 1026.5533, 1026.4719, 1026.3124, 1026.2006, 1026.0892, 1025.9348, 1025.7368, 1025.5707, 1025.4431, 1025.344, 1025.2213, 1025.1354, 1025.0767, 1024.9904, 1024.9012, 1024.8092, 1024.6816, 1024.2694, 1023.9551, 1023.9061, 1023.87744, 1023.85645, NaN, NaN, 1029.1758, 1029.1481, 1029.1133, 1029.0657, 1029.016, 1028.9684, 1028.9169, 1028.8668, 1028.8162, 1028.7618, 1028.7142, 1028.6687, 1028.6218, 1028.5748, 1028.5311, 1028.4807, 1028.4431, 1028.3931, 1028.3523, 1028.3019, 1028.2512, 1028.1951, 1028.152, 1028.1067, 1028.0614, 1028.0149, 1027.963, 1027.9095, 1027.854, 1027.8019, 1027.7494, 1027.694, 1027.6519, 1027.6078, 1027.5476, 1027.488, 1027.4271, 1027.3657, 1027.2979, 1027.244, 1027.1743, 1027.096, 1027.0326, 1026.9834, 1026.9174, 1026.8525, 1026.7694, 1026.6724, 1026.5773, 1026.5189, 1026.4073, 1026.2953, 1026.2002, 1026.012, 1025.8053, 1025.6649, 1025.567, 1025.4971, 1025.3615, 1025.2863, 1025.1816, 1025.1035, 1025.0612, 1024.9744, 1024.9038, 1024.8425, 1024.766, 1024.445, 1024.0774, 1023.9774, 1023.9327, 1023.9036, NaN, NaN, 1029.1805, 1029.1553, 1029.1173, 1029.069, 1029.0199, 1028.9607, 1028.9059, 1028.8479, 1028.791, 1028.7335, 1028.6744, 1028.6177, 1028.5646, 1028.5126, 1028.4591, 1028.4054, 1028.3455, 1028.2882, 1028.234, 1028.1793, 1028.1283, 1028.0758, 1028.0157, 1027.9574, 1027.8994, 1027.8347, 1027.787, 1027.7369, 1027.6823, 1027.6343, 1027.5793, 1027.5278, 1027.4651, 1027.3959, 1027.3438, 1027.2848, 1027.2097, 1027.1357, 1027.0872, 1027.0308, 1026.9509, 1026.8899, 1026.8169, 1026.7117, 1026.6201, 1026.5259, 1026.4625, 1026.3313, 1026.1969, 1025.9812, 1025.7748, 1025.6753, 1025.5076, 1025.418, 1025.3324, 1025.2681, 1025.1831, 1025.1208, 1025.0273, 1024.9358, 1024.8496, 1024.7957, 1024.6375, 1024.2732, 1024.1218, 1024.089, 1024.0626, 1024.0413, 1024.0255, NaN, NaN, 1029.1848, 1029.1586, 1029.1263, 1029.0797, 1029.033, 1028.9894, 1028.9386, 1028.8843, 1028.8232, 1028.7697, 1028.7166, 1028.6615, 1028.6094, 1028.5554, 1028.5059, 1028.4536, 1028.3972, 1028.339, 1028.2853, 1028.2313, 1028.1696, 1028.1077, 1028.0498, 1027.9966, 1027.9362, 1027.8861, 1027.8357, 1027.78, 1027.7263, 1027.6599, 1027.605, 1027.5557, 1027.4944, 1027.4288, 1027.3671, 1027.3079, 1027.2496, 1027.1743, 1027.0969, 1027.0222, 1026.9452, 1026.8601, 1026.797, 1026.6926, 1026.5703, 1026.455, 1026.3567, 1026.2714, 1026.1187, 1026.0065, 1025.7766, 1025.5859, 1025.4521, 1025.3501, 1025.2882, 1025.216, 1025.1306, 1025.0304, 1024.9199, 1024.7883, 1024.4597, 1024.2072, 1024.0574, 1024.0271, 1024.0, 1023.97797, 1023.9595, 1023.9478, NaN, NaN, 1029.1821, 1029.1494, 1029.114, 1029.0619, 1029.0035, 1028.951, 1028.893, 1028.8326, 1028.7716, 1028.7153, 1028.6611, 1028.6029, 1028.5459, 1028.4902, 1028.4369, 1028.3871, 1028.3323, 1028.2814, 1028.2322, 1028.1849, 1028.1299, 1028.0636, 1027.9972, 1027.9451, 1027.8967, 1027.8475, 1027.7969, 1027.7391, 1027.6813, 1027.6208, 1027.5647, 1027.5068, 1027.4462, 1027.3864, 1027.3365, 1027.2706, 1027.205, 1027.1428, 1027.0906, 1027.0243, 1026.9717, 1026.8892, 1026.8071, 1026.7275, 1026.6155, 1026.4857, 1026.3481, 1026.2236, 1026.1012, 1025.9678, 1025.7584, 1025.6193, 1025.5044, 1025.4159, 1025.3782, 1025.336, 1025.2253, 1025.1791, 1025.1307, 1025.0363, 1024.9379, 1024.8763, 1024.7485, 1024.4998, 1024.183, 1023.9789, 1023.9439, 1023.9219, 1023.9048, 1023.89136, 1023.87103, NaN, NaN, 1029.1858, 1029.1573, 1029.1213, 1029.0685, 1029.011, 1028.9476, 1028.895, 1028.8381, 1028.7864, 1028.7269, 1028.6664, 1028.6154, 1028.5627, 1028.5018, 1028.4465, 1028.3939, 1028.3472, 1028.2963, 1028.2389, 1028.18, 1028.1268, 1028.0781, 1028.029, 1027.9757, 1027.9241, 1027.8644, 1027.8102, 1027.7588, 1027.7083, 1027.6519, 1027.5975, 1027.5248, 1027.4562, 1027.397, 1027.3331, 1027.2743, 1027.205, 1027.1265, 1027.0599, 1026.9999, 1026.9211, 1026.8428, 1026.7756, 1026.6907, 1026.6147, 1026.5555, 1026.4056, 1026.2015, 1025.9674, 1025.8558, 1025.7576, 1025.6193, 1025.441, 1025.3905, 1025.335, 1025.2128, 1025.148, 1025.076, 1025.0066, 1024.9318, 1024.8145, 1024.4413, 1024.2046, 1023.99695, 1023.88434, 1023.8634, 1023.8428, 1023.82153, NaN, NaN, 1029.1948, 1029.166, 1029.1274, 1029.0748, 1029.0216, 1028.9712, 1028.9182, 1028.8636, 1028.8075, 1028.7511, 1028.6978, 1028.6467, 1028.5883, 1028.5283, 1028.4742, 1028.4222, 1028.3678, 1028.3112, 1028.2568, 1028.2, 1028.1472, 1028.0945, 1028.0369, 1027.9862, 1027.933, 1027.8815, 1027.8182, 1027.7584, 1027.7048, 1027.6467, 1027.5918, 1027.5367, 1027.4806, 1027.4279, 1027.364, 1027.2994, 1027.2196, 1027.1349, 1027.0757, 1027.0009, 1026.8961, 1026.8143, 1026.728, 1026.6462, 1026.5919, 1026.4554, 1026.2694, 1026.0674, 1025.9108, 1025.7495, 1025.5955, 1025.4999, 1025.4191, 1025.3711, 1025.2391, 1025.1768, 1025.0869, 1024.941, 1024.755, 1024.3647, 1024.2255, 1024.168, 1023.9261, 1023.8979, 1023.87946, 1023.8592, 1023.83356, 1023.8108, NaN, NaN, 1029.1675, 1029.1404, 1029.1057, 1029.0563, 1029.009, 1028.9551, 1028.9043, 1028.8574, 1028.8033, 1028.7555, 1028.7051, 1028.6572, 1028.6111, 1028.5543, 1028.5087, 1028.4622, 1028.4045, 1028.3447, 1028.2896, 1028.2406, 1028.1914, 1028.14, 1028.0898, 1028.0353, 1027.982, 1027.9286, 1027.8766, 1027.827, 1027.7761, 1027.7346, 1027.6748, 1027.6139, 1027.5706, 1027.5245, 1027.4678, 1027.4094, 1027.3501, 1027.294, 1027.2251, 1027.1544, 1027.0602, 1026.9844, 1026.9093, 1026.8153, 1026.7351, 1026.653, 1026.5546, 1026.458, 1026.3951, 1026.3022, 1026.1266, 1025.8882, 1025.7183, 1025.5677, 1025.4437, 1025.3804, 1025.2892, 1025.2438, 1025.2039, 1025.112, 1024.9886, 1024.8751, 1024.7819, 1024.5299, 1024.2328, 1024.1508, 1024.0128, 1023.9122, 1023.89624, 1023.8764, 1023.8522, 1023.82446, 1023.80707, NaN, NaN, 1029.1862, 1029.1577, 1029.1213, 1029.0662, 1029.0087, 1028.9565, 1028.903, 1028.8431, 1028.7948, 1028.7374, 1028.6874, 1028.6345, 1028.5844, 1028.5292, 1028.4723, 1028.4183, 1028.3611, 1028.3042, 1028.247, 1028.1869, 1028.1351, 1028.0839, 1028.0244, 1027.9806, 1027.9236, 1027.8613, 1027.8074, 1027.751, 1027.6958, 1027.633, 1027.5664, 1027.5089, 1027.4515, 1027.3881, 1027.3269, 1027.2561, 1027.1884, 1027.104, 1027.0259, 1026.897, 1026.817, 1026.7108, 1026.6183, 1026.5092, 1026.3898, 1026.241, 1026.0934, 1025.9578, 1025.7612, 1025.5919, 1025.451, 1025.2877, 1025.18, 1025.0975, 1024.9988, 1024.8987, 1024.7599, 1024.5753, 1024.2009, 1024.0054, 1023.9263, 1023.9017, 1023.8804, 1023.86084, 1023.8365, 1023.8162, NaN, NaN, 1029.1638, 1029.1355, 1029.0983, 1029.0469, 1028.9945, 1028.9388, 1028.8829, 1028.8317, 1028.7812, 1028.7324, 1028.6814, 1028.6278, 1028.5654, 1028.5167, 1028.4614, 1028.4126, 1028.3625, 1028.3141, 1028.2582, 1028.2034, 1028.1554, 1028.1055, 1028.0559, 1028.0011, 1027.953, 1027.9026, 1027.8441, 1027.7891, 1027.7338, 1027.6686, 1027.6138, 1027.5686, 1027.5195, 1027.4652, 1027.4034, 1027.34, 1027.2858, 1027.2297, 1027.1759, 1027.1055, 1027.041, 1026.939, 1026.8131, 1026.7075, 1026.6309, 1026.5183, 1026.4602, 1026.3019, 1026.1112, 1025.9744, 1025.8513, 1025.7029, 1025.5237, 1025.3385, 1025.1925, 1025.0951, 1024.9414, 1024.7386, 1024.4952, 1024.228, 1024.0293, 1023.96313, 1023.9395, 1023.9158, 1023.89435, 1023.86926, 1023.8471, 1023.82733, 1023.81024, NaN, NaN, 1029.1902, 1029.1611, 1029.1228, 1029.0737, 1029.0289, 1028.9749, 1028.9279, 1028.881, 1028.8293, 1028.777, 1028.7212, 1028.6656, 1028.614, 1028.5593, 1028.5105, 1028.457, 1028.4084, 1028.3527, 1028.3004, 1028.2468, 1028.1934, 1028.1489, 1028.1022, 1028.0461, 1027.9955, 1027.9426, 1027.8942, 1027.8438, 1027.7969, 1027.7421, 1027.6952, 1027.6469, 1027.6056, 1027.5464, 1027.4994, 1027.4542, 1027.3912, 1027.3367, 1027.2697, 1027.2057, 1027.1492, 1027.0782, 1027.0066, 1026.9103, 1026.7983, 1026.7008, 1026.6053, 1026.5238, 1026.4236, 1026.2891, 1026.1433, 1025.9758, 1025.837, 1025.6942, 1025.5471, 1025.4044, 1025.2699, 1025.164, 1025.0374, 1024.907, 1024.6117, 1024.3323, 1024.1156, 1024.0043, 1023.96454, 1023.94336, 1023.9226, 1023.905, 1023.88043, 1023.8523, 1023.8261, 1023.8115, NaN, NaN, 1029.1812, 1029.1514, 1029.1147, 1029.0685, 1029.0228, 1028.9728, 1028.9208, 1028.857, 1028.8026, 1028.7506, 1028.7006, 1028.6543, 1028.602, 1028.5466, 1028.4895, 1028.4403, 1028.3856, 1028.3297, 1028.271, 1028.2161, 1028.1682, 1028.1235, 1028.0723, 1028.0222, 1027.9695, 1027.9165, 1027.8705, 1027.8252, 1027.7776, 1027.723, 1027.6763, 1027.6271, 1027.5643, 1027.5114, 1027.4541, 1027.3896, 1027.3179, 1027.2499, 1027.2023, 1027.1411, 1027.0735, 1027.0027, 1026.9373, 1026.8657, 1026.7695, 1026.6735, 1026.6102, 1026.4425, 1026.3086, 1026.1672, 1026.0266, 1025.8534, 1025.6891, 1025.5658, 1025.4429, 1025.3059, 1025.1954, 1025.0071, 1024.8904, 1024.7971, 1024.5613, 1024.2981, 1024.1438, 1023.9922, 1023.95605, 1023.93176, 1023.9066, 1023.8817, 1023.8582, 1023.83905, 1023.82404, NaN, NaN, 1029.1747, 1029.1438, 1029.1088, 1029.0603, 1029.0145, 1028.9634, 1028.9164, 1028.868, 1028.8157, 1028.7656, 1028.7133, 1028.6611, 1028.6112, 1028.5619, 1028.5193, 1028.4694, 1028.4183, 1028.3661, 1028.3143, 1028.2539, 1028.2053, 1028.159, 1028.1135, 1028.0703, 1028.03, 1027.9797, 1027.9191, 1027.8667, 1027.8145, 1027.7594, 1027.7185, 1027.6609, 1027.6167, 1027.5625, 1027.4987, 1027.4375, 1027.3824, 1027.3098, 1027.2449, 1027.1903, 1027.1344, 1027.0798, 1027.011, 1026.9325, 1026.8448, 1026.7394, 1026.6619, 1026.5963, 1026.5177, 1026.4075, 1026.2728, 1026.112, 1025.9392, 1025.7723, 1025.6501, 1025.4929, 1025.3156, 1025.208, 1025.0868, 1024.9943, 1024.8965, 1024.762, 1024.5642, 1024.311, 1024.1206, 1023.96826, 1023.9488, 1023.92535, 1023.9047, 1023.8839, 1023.8574, 1023.83624, 1023.82166, NaN, NaN, 1029.1593, 1029.131, 1029.0953, 1029.0441, 1028.9888, 1028.9391, 1028.8876, 1028.8379, 1028.7869, 1028.7352, 1028.6838, 1028.632, 1028.583, 1028.5342, 1028.4878, 1028.4414, 1028.3905, 1028.3397, 1028.2959, 1028.2515, 1028.1969, 1028.1547, 1028.1086, 1028.0555, 1027.9983, 1027.9415, 1027.891, 1027.8416, 1027.7937, 1027.7428, 1027.695, 1027.6449, 1027.5884, 1027.5311, 1027.488, 1027.4336, 1027.378, 1027.3156, 1027.261, 1027.2025, 1027.1448, 1027.082, 1027.0139, 1026.9434, 1026.8927, 1026.836, 1026.7661, 1026.6956, 1026.6207, 1026.5261, 1026.4407, 1026.3022, 1026.0876, 1025.9001, 1025.7373, 1025.5935, 1025.3889, 1025.2887, 1025.1351, 1025.0038, 1024.8717, 1024.7676, 1024.5149, 1024.2118, 1024.0084, 1023.9721, 1023.9491, 1023.9285, 1023.9047, 1023.8798, 1023.8535, 1023.82825, 1023.81396, NaN, NaN, 1029.159, 1029.1261, 1029.0863, 1029.0332, 1028.9812, 1028.9276, 1028.8707, 1028.8193, 1028.7692, 1028.7108, 1028.6548, 1028.5975, 1028.5459, 1028.4878, 1028.4279, 1028.3812, 1028.3326, 1028.2819, 1028.2223, 1028.1613, 1028.0978, 1028.0361, 1027.9728, 1027.9193, 1027.863, 1027.8109, 1027.7559, 1027.6981, 1027.646, 1027.5868, 1027.5209, 1027.443, 1027.374, 1027.3215, 1027.2695, 1027.2142, 1027.151, 1027.0868, 1027.028, 1026.978, 1026.9215, 1026.8483, 1026.7742, 1026.7119, 1026.6234, 1026.5222, 1026.3927, 1026.1924, 1025.9541, 1025.8302, 1025.7118, 1025.6277, 1025.4678, 1025.3629, 1025.2731, 1025.1104, 1024.9867, 1024.8169, 1024.6573, 1024.3685, 1024.0446, 1023.9596, 1023.9318, 1023.90735, 1023.88513, 1023.86646, 1023.8388, 1023.8236, NaN, NaN, 1029.1371, 1029.111, 1029.077, 1029.024, 1028.968, 1028.9167, 1028.8645, 1028.7986, 1028.7456, 1028.6938, 1028.6426, 1028.5842, 1028.537, 1028.4727, 1028.4246, 1028.3707, 1028.3271, 1028.274, 1028.2163, 1028.1534, 1028.0953, 1028.0433, 1027.9822, 1027.9171, 1027.864, 1027.8121, 1027.7635, 1027.7141, 1027.6586, 1027.6044, 1027.5476, 1027.4843, 1027.4281, 1027.362, 1027.3007, 1027.2554, 1027.2091, 1027.1415, 1027.0764, 1027.0182, 1026.9629, 1026.901, 1026.8351, 1026.7534, 1026.6866, 1026.5782, 1026.4116, 1026.2687, 1026.1775, 1026.0608, 1025.8867, 1025.7188, 1025.6023, 1025.477, 1025.3478, 1025.2068, 1025.1117, 1025.0006, 1024.7893, 1024.591, 1024.3289, 1024.0027, 1023.9571, 1023.93225, 1023.9074, 1023.883, 1023.8678, 1023.84827, NaN, NaN, 1029.1714, 1029.1389, 1029.0961, 1029.038, 1028.9946, 1028.9481, 1028.8972, 1028.8398, 1028.7843, 1028.7279, 1028.6753, 1028.6188, 1028.5688, 1028.5161, 1028.4602, 1028.399, 1028.3503, 1028.2999, 1028.2451, 1028.1926, 1028.1333, 1028.0768, 1028.0215, 1027.9662, 1027.9114, 1027.8541, 1027.8055, 1027.7599, 1027.7108, 1027.6564, 1027.5988, 1027.5377, 1027.4756, 1027.415, 1027.3519, 1027.2893, 1027.2358, 1027.1799, 1027.122, 1027.0516, 1026.9823, 1026.9116, 1026.8466, 1026.7823, 1026.7211, 1026.6663, 1026.559, 1026.4015, 1026.2229, 1026.0459, 1025.8892, 1025.696, 1025.5189, 1025.3823, 1025.2083, 1025.0931, 1024.9626, 1024.823, 1024.6703, 1024.5255, 1024.208, 1024.0583, 1024.0374, 1024.0099, 1023.98517, 1023.9631, 1023.94086, 1023.9296, NaN, NaN, 1029.1836, 1029.1558, 1029.1136, 1029.0543, 1028.9955, 1028.948, 1028.9005, 1028.852, 1028.8014, 1028.7518, 1028.6954, 1028.6406, 1028.586, 1028.534, 1028.4664, 1028.4199, 1028.3743, 1028.3237, 1028.2745, 1028.2225, 1028.1666, 1028.1023, 1028.0475, 1027.9998, 1027.947, 1027.8889, 1027.8461, 1027.7942, 1027.7423, 1027.6909, 1027.6401, 1027.5775, 1027.5206, 1027.4705, 1027.4019, 1027.3458, 1027.2998, 1027.2382, 1027.167, 1027.1011, 1027.0297, 1026.9583, 1026.9003, 1026.8468, 1026.7988, 1026.7433, 1026.6813, 1026.6152, 1026.5299, 1026.3555, 1026.1882, 1025.9862, 1025.7817, 1025.5675, 1025.4209, 1025.2722, 1025.1736, 1025.0521, 1024.9094, 1024.7488, 1024.6533, 1024.5576, 1024.3197, 1024.1034, 1023.99316, 1023.9684, 1023.9484, 1023.92035, 1023.90393, NaN, NaN, 1029.1731, 1029.1462, 1029.102, 1029.048, 1028.9954, 1028.9409, 1028.8895, 1028.8362, 1028.7856, 1028.7313, 1028.6776, 1028.6267, 1028.5717, 1028.5138, 1028.4506, 1028.4033, 1028.3542, 1028.3015, 1028.2395, 1028.1805, 1028.1195, 1028.0634, 1028.0099, 1027.9557, 1027.907, 1027.8544, 1027.7999, 1027.7426, 1027.6887, 1027.6266, 1027.5808, 1027.5204, 1027.457, 1027.3997, 1027.361, 1027.316, 1027.2549, 1027.201, 1027.134, 1027.0681, 1027.0032, 1026.9427, 1026.8887, 1026.8381, 1026.7853, 1026.72, 1026.6536, 1026.543, 1026.3939, 1026.2443, 1026.0593, 1025.9247, 1025.764, 1025.6305, 1025.5178, 1025.3815, 1025.2657, 1025.1974, 1025.1222, 1024.9767, 1024.8376, 1024.7291, 1024.5986, 1024.4716, 1024.3936, 1024.2397, 1024.058, 1024.0283, 1023.99493, 1023.9702, 1023.9512, NaN, NaN, 1029.1759, 1029.1481, 1029.1128, 1029.0605, 1029.0045, 1028.9513, 1028.8955, 1028.8472, 1028.8046, 1028.7516, 1028.702, 1028.655, 1028.5936, 1028.5371, 1028.4747, 1028.4054, 1028.3513, 1028.2933, 1028.2341, 1028.1885, 1028.14, 1028.0881, 1028.0325, 1027.9769, 1027.9141, 1027.8588, 1027.8036, 1027.7511, 1027.7013, 1027.6426, 1027.5856, 1027.5264, 1027.4674, 1027.3998, 1027.3419, 1027.2906, 1027.2299, 1027.16, 1027.0939, 1027.0283, 1026.9617, 1026.907, 1026.8556, 1026.802, 1026.7432, 1026.6777, 1026.606, 1026.4799, 1026.339, 1026.2015, 1026.036, 1025.8806, 1025.7302, 1025.5747, 1025.4062, 1025.285, 1025.1787, 1025.0883, 1024.9268, 1024.7795, 1024.6182, 1024.503, 1024.4182, 1024.1951, 1024.0236, 1023.9866, 1023.95844, 1023.9405, NaN, NaN, 1029.1825, 1029.1509, 1029.1149, 1029.0629, 1029.0045, 1028.9451, 1028.8911, 1028.8317, 1028.7743, 1028.7228, 1028.6632, 1028.6147, 1028.5698, 1028.516, 1028.462, 1028.407, 1028.3542, 1028.3053, 1028.2546, 1028.2087, 1028.1611, 1028.114, 1028.0559, 1028.0021, 1027.9531, 1027.896, 1027.8439, 1027.7886, 1027.7347, 1027.6877, 1027.6387, 1027.5874, 1027.5267, 1027.4637, 1027.4005, 1027.3584, 1027.3154, 1027.267, 1027.1973, 1027.1217, 1027.0497, 1026.995, 1026.9349, 1026.867, 1026.8046, 1026.7401, 1026.656, 1026.5741, 1026.4542, 1026.3015, 1026.1902, 1026.0219, 1025.8519, 1025.7457, 1025.6329, 1025.5048, 1025.3184, 1025.178, 1025.043, 1024.9073, 1024.7993, 1024.6747, 1024.5739, 1024.441, 1024.2689, 1024.0455, 1024.0138, 1023.99066, 1023.9644, 1023.94684, NaN, NaN, 1029.1604, 1029.1326, 1029.091, 1029.0378, 1028.9882, 1028.9314, 1028.8657, 1028.8058, 1028.7484, 1028.6954, 1028.6383, 1028.5835, 1028.5239, 1028.4645, 1028.4062, 1028.3402, 1028.2755, 1028.212, 1028.1564, 1028.1079, 1028.061, 1028.0132, 1027.9498, 1027.8937, 1027.8376, 1027.781, 1027.7216, 1027.6532, 1027.5986, 1027.5339, 1027.4624, 1027.4008, 1027.3386, 1027.2798, 1027.2336, 1027.1729, 1027.1019, 1027.0233, 1026.9672, 1026.8888, 1026.8345, 1026.7563, 1026.6697, 1026.5709, 1026.4443, 1026.3246, 1026.1753, 1026.0184, 1025.879, 1025.6669, 1025.4832, 1025.3357, 1025.2207, 1025.1044, 1025.0023, 1024.9131, 1024.7571, 1024.6635, 1024.5411, 1024.4181, 1024.1974, 1024.0804, 1024.0559, 1024.035, 1024.0161, 1023.98987, 1023.97064, NaN, NaN, 1029.188, 1029.1615, 1029.123, 1029.0707, 1029.0215, 1028.9698, 1028.918, 1028.8657, 1028.814, 1028.7615, 1028.7047, 1028.6465, 1028.5948, 1028.5375, 1028.4801, 1028.4236, 1028.3668, 1028.3108, 1028.253, 1028.1915, 1028.1381, 1028.0851, 1028.0331, 1027.9827, 1027.9285, 1027.8749, 1027.8214, 1027.7714, 1027.7135, 1027.653, 1027.5984, 1027.5464, 1027.4911, 1027.4349, 1027.3798, 1027.3098, 1027.2406, 1027.1884, 1027.1222, 1027.0693, 1027.0184, 1026.9578, 1026.9069, 1026.8369, 1026.7656, 1026.6857, 1026.5956, 1026.4814, 1026.3639, 1026.263, 1026.0757, 1025.9543, 1025.7444, 1025.5826, 1025.4564, 1025.359, 1025.2089, 1025.1049, 1024.9454, 1024.7924, 1024.6616, 1024.5201, 1024.4451, 1024.2979, 1024.1198, 1024.0754, 1024.0515, 1024.032, 1024.0106, 1023.986, NaN, NaN, 1029.2056, 1029.1726, 1029.1321, 1029.0793, 1029.0192, 1028.9631, 1028.9062, 1028.8542, 1028.8013, 1028.7496, 1028.6981, 1028.6461, 1028.595, 1028.5399, 1028.4784, 1028.4246, 1028.3636, 1028.3114, 1028.257, 1028.1968, 1028.149, 1028.095, 1028.0413, 1027.9828, 1027.9247, 1027.8691, 1027.8184, 1027.7631, 1027.7002, 1027.6339, 1027.5648, 1027.4984, 1027.4387, 1027.3729, 1027.301, 1027.229, 1027.1539, 1027.0767, 1027.001, 1026.9393, 1026.8689, 1026.7963, 1026.7273, 1026.6482, 1026.5535, 1026.4492, 1026.3112, 1026.1482, 1025.9958, 1025.87, 1025.7032, 1025.6229, 1025.5226, 1025.4124, 1025.309, 1025.2014, 1025.1244, 1025.0151, 1024.831, 1024.7183, 1024.6432, 1024.5609, 1024.4564, 1024.2938, 1024.1024, 1024.0723, 1024.0459, 1024.0248, 1024.0123, NaN, NaN, 1029.1824, 1029.1532, 1029.1149, 1029.069, 1029.0289, 1028.9807, 1028.935, 1028.887, 1028.8392, 1028.7882, 1028.7339, 1028.6891, 1028.6416, 1028.5895, 1028.5372, 1028.4893, 1028.4387, 1028.3883, 1028.3401, 1028.2903, 1028.2407, 1028.1891, 1028.1372, 1028.0862, 1028.027, 1027.9719, 1027.918, 1027.8624, 1027.8201, 1027.7698, 1027.7218, 1027.6722, 1027.6183, 1027.5647, 1027.5042, 1027.4469, 1027.3888, 1027.3246, 1027.2627, 1027.1951, 1027.1185, 1027.0518, 1026.9684, 1026.8843, 1026.8002, 1026.7164, 1026.6168, 1026.5316, 1026.3953, 1026.2765, 1026.1641, 1026.0345, 1025.8661, 1025.6985, 1025.5651, 1025.4205, 1025.3138, 1025.2013, 1025.0809, 1024.9442, 1024.8096, 1024.6882, 1024.5729, 1024.4539, 1024.183, 1024.1042, 1024.0608, 1024.0361, 1024.0112, 1023.33923, 1022.77374, 1022.87177, NaN, NaN, 1027.1027, 1027.0527, 1026.9895, 1026.8816, 1026.8083, 1026.7448, 1026.6655, 1026.5532, 1026.4542, 1026.4225, 1026.3198, 1026.0619, 1026.3538, 1026.2589, 1026.2379, 1026.1927, 1026.0197, 1026.5497, 1028.2483, 1028.1919, 1028.1349, 1028.0778, 1028.0194, 1027.9597, 1027.895, 1027.8373, 1027.79, 1027.7281, 1027.6746, 1027.6151, 1027.5662, 1027.5098, 1027.4513, 1027.3838, 1027.325, 1027.2604, 1027.1897, 1027.111, 1027.0371, 1026.9642, 1026.8978, 1026.8147, 1026.7201, 1026.6237, 1026.4954, 1026.287, 1026.1293, 1026.0052, 1025.8566, 1025.7249, 1025.5902, 1025.4452, 1025.3221, 1025.1984, 1025.083, 1024.9622, 1024.7975, 1024.6351, 1024.537, 1024.2335, 1024.1045, 1024.0698, 1024.0321, 1023.99316, 1023.918, 1023.87006, 1023.85315, NaN, NaN, 1029.1819, 1029.1543, 1029.1207, 1029.0773, 1029.0374, 1028.9895, 1028.938, 1028.8892, 1028.8445, 1028.7977, 1028.7533, 1028.7012, 1028.6469, 1028.5953, 1028.5454, 1028.4901, 1028.4358, 1028.3768, 1028.3225, 1028.2682, 1028.2158, 1028.1595, 1028.102, 1028.0414, 1027.9855, 1027.9337, 1027.8846, 1027.8323, 1027.774, 1027.7223, 1027.6632, 1027.6145, 1027.5653, 1027.5105, 1027.4536, 1027.3982, 1027.3367, 1027.2698, 1027.2148, 1027.1434, 1027.0583, 1026.9688, 1026.8986, 1026.8114, 1026.7194, 1026.6346, 1026.5344, 1026.4172, 1026.2883, 1026.1625, 1026.0048, 1025.8265, 1025.6823, 1025.5494, 1025.4243, 1025.2777, 1025.1685, 1025.0848, 1024.9729, 1024.8093, 1024.6874, 1024.5876, 1024.4196, 1024.1211, 1024.0579, 1024.0299, 1023.9956, 1023.9496, 1023.8636, 1023.8369, NaN, NaN, 1029.2056, 1029.1698, 1029.1311, 1029.0841, 1029.034, 1028.9757, 1028.9218, 1028.8751, 1028.8229, 1028.765, 1028.7142, 1028.6672, 1028.6173, 1028.5658, 1028.5121, 1028.4548, 1028.3873, 1028.3318, 1028.2836, 1028.2334, 1028.186, 1028.1364, 1028.0844, 1028.0265, 1027.9681, 1027.9054, 1027.8444, 1027.7909, 1027.7362, 1027.6774, 1027.616, 1027.5663, 1027.5187, 1027.4633, 1027.3944, 1027.3296, 1027.2681, 1027.2109, 1027.151, 1027.0874, 1027.0145, 1026.9387, 1026.8582, 1026.7465, 1026.6467, 1026.5366, 1026.3909, 1026.2695, 1026.1509, 1026.0287, 1025.8768, 1025.6686, 1025.4951, 1025.3572, 1025.255, 1025.1534, 1025.062, 1024.9601, 1024.8486, 1024.718, 1024.561, 1024.3793, 1024.1031, 1024.0652, 1024.0062, 1023.9654, 1023.87146, 1023.76965, 1023.7216, 1023.7038, NaN, NaN, 1029.1951, 1029.1686, 1029.1338, 1029.084, 1029.0255, 1028.9711, 1028.9149, 1028.8619, 1028.8079, 1028.7574, 1028.706, 1028.6536, 1028.6033, 1028.5447, 1028.4911, 1028.4344, 1028.384, 1028.3314, 1028.2836, 1028.2255, 1028.1709, 1028.1116, 1028.0555, 1027.9834, 1027.9183, 1027.859, 1027.8048, 1027.7446, 1027.6831, 1027.6194, 1027.5607, 1027.5001, 1027.45, 1027.3882, 1027.3225, 1027.2614, 1027.1863, 1027.1002, 1027.0404, 1026.9794, 1026.9146, 1026.8278, 1026.7101, 1026.5908, 1026.4713, 1026.3269, 1026.1584, 1026.0688, 1025.8171, 1025.6188, 1025.4681, 1025.3152, 1025.1962, 1025.0707, 1024.9707, 1024.8568, 1024.716, 1024.5524, 1024.2819, 1024.0677, 1024.0024, 1023.91315, 1023.85223, 1023.7871, 1023.7425, 1023.70294, 1023.6669, NaN, NaN, 1029.2183, 1029.1901, 1029.1539, 1029.1084, 1029.0638, 1029.0116, 1028.9596, 1028.9114, 1028.858, 1028.8073, 1028.7563, 1028.7057, 1028.6564, 1028.6085, 1028.5544, 1028.5062, 1028.4521, 1028.3926, 1028.3458, 1028.2966, 1028.2467, 1028.199, 1028.1526, 1028.1052, 1028.0509, 1027.9956, 1027.9368, 1027.8784, 1027.8243, 1027.7795, 1027.7284, 1027.6572, 1027.5887, 1027.5345, 1027.4811, 1027.4288, 1027.3741, 1027.3235, 1027.2705, 1027.2048, 1027.134, 1027.0597, 1026.9883, 1026.9156, 1026.8177, 1026.7164, 1026.632, 1026.5442, 1026.4297, 1026.3182, 1026.2056, 1026.0596, 1025.9408, 1025.6888, 1025.5078, 1025.3514, 1025.2622, 1025.1376, 1025.0498, 1024.948, 1024.794, 1024.5989, 1024.3362, 1024.0897, 1024.0116, 1023.9668, 1023.94556, 1023.90814, 1023.8532, 1023.7462, 1023.69745, NaN, NaN, 1029.1979, 1029.1714, 1029.1365, 1029.0914, 1029.0492, 1029.0062, 1028.9557, 1028.9132, 1028.8625, 1028.809, 1028.7599, 1028.7117, 1028.6705, 1028.627, 1028.5742, 1028.5288, 1028.4797, 1028.4315, 1028.3851, 1028.3367, 1028.2853, 1028.2397, 1028.1946, 1028.1538, 1028.1062, 1028.0554, 1027.9978, 1027.9537, 1027.8994, 1027.8463, 1027.7933, 1027.7396, 1027.6923, 1027.6405, 1027.583, 1027.5208, 1027.469, 1027.4146, 1027.353, 1027.2911, 1027.2324, 1027.1733, 1027.113, 1027.0535, 1026.9913, 1026.929, 1026.8536, 1026.7533, 1026.6653, 1026.5682, 1026.4741, 1026.3558, 1026.2263, 1026.1129, 1026.0022, 1025.9304, 1025.8315, 1025.6974, 1025.5515, 1025.4197, 1025.3068, 1025.1886, 1025.0574, 1024.9268, 1024.8187, 1024.6147, 1024.3414, 1024.0525, 1023.9776, 1023.9523, 1023.92487, 1023.89343, 1023.8251, NaN, NaN, 1029.2056, 1029.1742, 1029.1393, 1029.0859, 1029.0317, 1028.9747, 1028.9204, 1028.8667, 1028.8103, 1028.7559, 1028.6996, 1028.6473, 1028.593, 1028.5374, 1028.4802, 1028.4243, 1028.37, 1028.318, 1028.266, 1028.2146, 1028.1649, 1028.1084, 1028.0559, 1028.0072, 1027.9619, 1027.9113, 1027.8599, 1027.7998, 1027.7404, 1027.688, 1027.6437, 1027.5951, 1027.5249, 1027.4681, 1027.4132, 1027.3536, 1027.3026, 1027.2546, 1027.1908, 1027.1161, 1027.0364, 1026.9498, 1026.867, 1026.772, 1026.6616, 1026.5334, 1026.4338, 1026.3196, 1026.2236, 1026.1035, 1025.9862, 1025.8441, 1025.7045, 1025.5632, 1025.4058, 1025.3165, 1025.201, 1025.0951, 1024.9543, 1024.8737, 1024.7563, 1024.5712, 1024.3878, 1024.065, 1024.0044, 1023.9719, 1023.94025, 1023.90027, 1023.8211, 1023.7925, NaN, NaN, 1029.2107, 1029.1825, 1029.1456, 1029.0908, 1029.0342, 1028.9812, 1028.9293, 1028.8787, 1028.8252, 1028.7767, 1028.7279, 1028.6759, 1028.6249, 1028.5767, 1028.5239, 1028.4719, 1028.4236, 1028.3696, 1028.3108, 1028.2592, 1028.1973, 1028.1422, 1028.089, 1028.0295, 1027.975, 1027.9126, 1027.8505, 1027.7845, 1027.7087, 1027.6478, 1027.5828, 1027.5062, 1027.4321, 1027.3774, 1027.3102, 1027.2441, 1027.1736, 1027.1053, 1027.0331, 1026.9603, 1026.8815, 1026.8087, 1026.696, 1026.5579, 1026.4458, 1026.2793, 1026.1268, 1025.9608, 1025.8234, 1025.6335, 1025.4741, 1025.3484, 1025.255, 1025.1116, 1024.9703, 1024.8705, 1024.78, 1024.5677, 1024.428, 1024.3308, 1024.1941, 1024.1184, 1024.0305, 1023.92395, 1023.8574, 1023.8284, 1023.81354, NaN, NaN, 1029.2263, 1029.1989, 1029.1608, 1029.1104, 1029.0594, 1029.0042, 1028.9478, 1028.8899, 1028.8392, 1028.7836, 1028.7269, 1028.6747, 1028.6241, 1028.5739, 1028.517, 1028.4675, 1028.4161, 1028.365, 1028.3143, 1028.2607, 1028.2036, 1028.1466, 1028.0956, 1028.0438, 1027.9943, 1027.9419, 1027.8855, 1027.8328, 1027.7831, 1027.7205, 1027.6604, 1027.6118, 1027.5619, 1027.5023, 1027.4459, 1027.3777, 1027.3171, 1027.2496, 1027.1898, 1027.1165, 1027.0404, 1026.9624, 1026.8827, 1026.786, 1026.6906, 1026.5563, 1026.3823, 1026.1809, 1026.0239, 1025.8798, 1025.7681, 1025.6389, 1025.5059, 1025.3774, 1025.2712, 1025.156, 1025.0128, 1024.9073, 1024.7926, 1024.6017, 1024.4636, 1024.3448, 1024.2166, 1024.0723, 1024.0038, 1023.96277, 1023.91876, 1023.8949, NaN, NaN, 1029.2084, 1029.178, 1029.1422, 1029.09, 1029.0332, 1028.9755, 1028.9247, 1028.8672, 1028.8098, 1028.7567, 1028.7013, 1028.6454, 1028.5933, 1028.544, 1028.4922, 1028.4386, 1028.3895, 1028.3383, 1028.2869, 1028.2349, 1028.1881, 1028.139, 1028.0853, 1028.0333, 1027.9761, 1027.9083, 1027.8602, 1027.8088, 1027.7542, 1027.6927, 1027.6393, 1027.581, 1027.5237, 1027.4652, 1027.402, 1027.3381, 1027.2797, 1027.1953, 1027.1194, 1027.0626, 1026.9966, 1026.921, 1026.8406, 1026.752, 1026.6407, 1026.5421, 1026.3978, 1026.2273, 1026.0791, 1025.928, 1025.7864, 1025.6555, 1025.564, 1025.4584, 1025.3256, 1025.2289, 1025.141, 1025.0697, 1024.9724, 1024.8483, 1024.683, 1024.6154, 1024.4935, 1024.31, 1024.1628, 1024.0841, 1023.9737, 1023.92755, 1023.8968, NaN, NaN, 1029.2197, 1029.1919, 1029.1571, 1029.1085, 1029.0615, 1029.0137, 1028.9609, 1028.9119, 1028.8615, 1028.8104, 1028.7607, 1028.712, 1028.6602, 1028.6062, 1028.5527, 1028.4995, 1028.4475, 1028.3938, 1028.3397, 1028.2899, 1028.2401, 1028.1837, 1028.1327, 1028.0789, 1028.0189, 1027.9559, 1027.9095, 1027.8551, 1027.8005, 1027.7511, 1027.6978, 1027.6477, 1027.5968, 1027.5488, 1027.508, 1027.4517, 1027.4075, 1027.3417, 1027.2758, 1027.2189, 1027.1566, 1027.0859, 1027.038, 1026.9708, 1026.9147, 1026.8014, 1026.6995, 1026.5732, 1026.4589, 1026.3197, 1026.1748, 1026.0334, 1025.9116, 1025.779, 1025.6469, 1025.5505, 1025.4602, 1025.3309, 1025.235, 1025.1748, 1025.0845, 1024.9647, 1024.8716, 1024.7539, 1024.6245, 1024.5116, 1024.3785, 1024.1409, 1023.9984, 1023.9596, 1023.9343, 1023.91833, NaN, NaN, 1029.2227, 1029.1931, 1029.152, 1029.1008, 1029.0542, 1029.0039, 1028.9434, 1028.8835, 1028.8262, 1028.7737, 1028.7195, 1028.6617, 1028.6053, 1028.5463, 1028.4886, 1028.428, 1028.3755, 1028.3228, 1028.2747, 1028.2197, 1028.1692, 1028.1193, 1028.0651, 1028.0183, 1027.9626, 1027.9158, 1027.8651, 1027.8063, 1027.7502, 1027.6962, 1027.6409, 1027.5836, 1027.5298, 1027.467, 1027.3909, 1027.3342, 1027.2731, 1027.2091, 1027.146, 1027.0762, 1027.0048, 1026.9347, 1026.833, 1026.7405, 1026.6241, 1026.5162, 1026.3948, 1026.2491, 1026.1381, 1025.9296, 1025.7224, 1025.6196, 1025.4938, 1025.4197, 1025.3538, 1025.2363, 1025.1388, 1025.0667, 1024.9775, 1024.8593, 1024.7313, 1024.5498, 1024.4442, 1024.2716, 1024.0798, 1024.0043, 1023.96027, 1023.9362, 1023.911, 1023.8951, NaN, NaN, 1029.2385, 1029.2089, 1029.1733, 1029.1277, 1029.0776, 1029.028, 1028.9784, 1028.93, 1028.8794, 1028.8315, 1028.7839, 1028.7307, 1028.6754, 1028.6248, 1028.5715, 1028.5227, 1028.4698, 1028.4155, 1028.3661, 1028.3159, 1028.2601, 1028.2039, 1028.1484, 1028.0868, 1028.0288, 1027.9717, 1027.909, 1027.8524, 1027.8, 1027.7494, 1027.6897, 1027.637, 1027.5771, 1027.5186, 1027.4675, 1027.4135, 1027.353, 1027.2964, 1027.2413, 1027.1829, 1027.1149, 1027.0338, 1026.9543, 1026.8577, 1026.766, 1026.6893, 1026.5865, 1026.4818, 1026.3145, 1026.1715, 1026.0026, 1025.8903, 1025.7388, 1025.5305, 1025.3928, 1025.2631, 1025.1276, 1025.04, 1024.9138, 1024.7927, 1024.6299, 1024.4224, 1024.218, 1024.0759, 1024.0306, 1024.0013, 1023.9687, 1023.92957, 1023.8957, 1023.8821, NaN, NaN, 1029.2394, 1029.2128, 1029.1753, 1029.1293, 1029.0798, 1029.0306, 1028.9728, 1028.9232, 1028.8695, 1028.817, 1028.7623, 1028.7019, 1028.6409, 1028.582, 1028.5295, 1028.4779, 1028.426, 1028.369, 1028.3099, 1028.2556, 1028.2025, 1028.145, 1028.0924, 1028.0372, 1027.9794, 1027.9216, 1027.8645, 1027.8064, 1027.7513, 1027.6945, 1027.6312, 1027.5757, 1027.5223, 1027.4672, 1027.4062, 1027.3353, 1027.271, 1027.1997, 1027.1212, 1027.0383, 1026.9407, 1026.8539, 1026.7537, 1026.6069, 1026.4542, 1026.2913, 1026.1257, 1026.0177, 1025.937, 1025.8104, 1025.6943, 1025.5299, 1025.4039, 1025.2909, 1025.1569, 1025.058, 1024.9913, 1024.8665, 1024.6887, 1024.436, 1024.2517, 1024.111, 1024.0791, 1024.0537, 1024.0128, 1023.93823, 1023.88947, 1023.8679, NaN, NaN, 1029.2421, 1029.2164, 1029.1807, 1029.1372, 1029.0892, 1029.0392, 1028.9917, 1028.947, 1028.8966, 1028.8464, 1028.7972, 1028.7483, 1028.6998, 1028.6511, 1028.6, 1028.5474, 1028.498, 1028.4481, 1028.3988, 1028.3461, 1028.2909, 1028.2328, 1028.1782, 1028.1293, 1028.0834, 1028.0265, 1027.9724, 1027.9192, 1027.8584, 1027.8054, 1027.7513, 1027.6925, 1027.6335, 1027.577, 1027.5226, 1027.4633, 1027.4031, 1027.3336, 1027.2688, 1027.1926, 1027.132, 1027.0642, 1026.9625, 1026.8429, 1026.7554, 1026.6492, 1026.5278, 1026.4001, 1026.26, 1026.0887, 1025.908, 1025.7493, 1025.6193, 1025.4718, 1025.3197, 1025.232, 1025.1063, 1025.0238, 1024.9666, 1024.8854, 1024.7799, 1024.6484, 1024.4669, 1024.2339, 1024.096, 1024.0717, 1024.0305, 1023.93994, 1023.9061, 1023.872, 1023.8493, NaN, NaN, 1029.2366, 1029.2074, 1029.173, 1029.1285, 1029.0841, 1029.0391, 1028.9937, 1028.9489, 1028.9038, 1028.8588, 1028.8058, 1028.7556, 1028.6989, 1028.6469, 1028.5933, 1028.5443, 1028.493, 1028.4393, 1028.3804, 1028.3247, 1028.2789, 1028.2285, 1028.1742, 1028.122, 1028.069, 1028.015, 1027.9519, 1027.8964, 1027.8464, 1027.8024, 1027.755, 1027.7067, 1027.6573, 1027.6, 1027.5408, 1027.4916, 1027.4342, 1027.3773, 1027.3236, 1027.2712, 1027.2139, 1027.1366, 1027.066, 1026.9698, 1026.877, 1026.7637, 1026.6514, 1026.5308, 1026.3828, 1026.2562, 1026.1152, 1025.9207, 1025.777, 1025.6442, 1025.5336, 1025.4059, 1025.2766, 1025.1753, 1025.0963, 1024.9724, 1024.8733, 1024.7347, 1024.5674, 1024.4504, 1024.1471, 1024.0427, 1023.9731, 1023.91455, 1023.88544, 1023.86395, 1023.84906, NaN, NaN, 1029.2422, 1029.2156, 1029.1833, 1029.1355, 1029.082, 1029.0295, 1028.9769, 1028.9246, 1028.8723, 1028.8239, 1028.7731, 1028.7222, 1028.6747, 1028.6179, 1028.563, 1028.5112, 1028.4553, 1028.3953, 1028.3376, 1028.2809, 1028.2233, 1028.1707, 1028.119, 1028.0642, 1028.0021, 1027.9453, 1027.8893, 1027.8373, 1027.786, 1027.7303, 1027.6735, 1027.6119, 1027.5526, 1027.4939, 1027.4308, 1027.3694, 1027.2961, 1027.2216, 1027.1348, 1027.0791, 1027.0072, 1026.9348, 1026.8539, 1026.773, 1026.6891, 1026.542, 1026.3826, 1026.2354, 1026.0532, 1025.8798, 1025.705, 1025.5583, 1025.4487, 1025.3931, 1025.2083, 1025.0734, 1024.9546, 1024.8617, 1024.6664, 1024.5437, 1024.4247, 1024.2128, 1024.0768, 1024.025, 1023.9491, 1023.8948, 1023.85693, 1023.8367, NaN, NaN, 1029.2471, 1029.2184, 1029.1838, 1029.1411, 1029.0956, 1029.0447, 1028.9924, 1028.9462, 1028.8982, 1028.8485, 1028.8026, 1028.7552, 1028.7057, 1028.6576, 1028.613, 1028.5637, 1028.5095, 1028.4602, 1028.4141, 1028.3616, 1028.3137, 1028.2653, 1028.2137, 1028.1688, 1028.1224, 1028.0742, 1028.0178, 1027.9626, 1027.9125, 1027.8633, 1027.81, 1027.7537, 1027.7026, 1027.6462, 1027.5956, 1027.5385, 1027.479, 1027.4188, 1027.3656, 1027.3119, 1027.2395, 1027.1495, 1027.0759, 1026.9857, 1026.8704, 1026.7511, 1026.6014, 1026.4717, 1026.3346, 1026.2308, 1025.9573, 1025.8408, 1025.6741, 1025.5277, 1025.4159, 1025.3169, 1025.182, 1025.0571, 1024.9174, 1024.7596, 1024.6421, 1024.4846, 1024.3313, 1024.2556, 1024.1239, 1024.0643, 1024.0206, 1023.921, 1023.8776, 1023.8487, 1023.8252, NaN, NaN, 1029.2434, 1029.2153, 1029.1791, 1029.1305, 1029.0757, 1029.0247, 1028.9714, 1028.9209, 1028.8695, 1028.8198, 1028.7693, 1028.7177, 1028.6628, 1028.6091, 1028.5532, 1028.5033, 1028.4506, 1028.4009, 1028.3496, 1028.2944, 1028.2405, 1028.1832, 1028.1255, 1028.072, 1028.0217, 1027.9603, 1027.9048, 1027.8536, 1027.7959, 1027.7393, 1027.6906, 1027.6399, 1027.5876, 1027.5353, 1027.4736, 1027.4178, 1027.3561, 1027.2837, 1027.2094, 1027.1387, 1027.0623, 1026.9734, 1026.8806, 1026.7953, 1026.7084, 1026.617, 1026.4207, 1026.2529, 1026.1119, 1026.0006, 1025.8633, 1025.7036, 1025.577, 1025.4172, 1025.2802, 1025.1564, 1025.063, 1024.9073, 1024.7684, 1024.6135, 1024.4559, 1024.27, 1024.0892, 1024.0509, 1023.9854, 1023.89923, 1023.8496, 1023.81573, 1023.7918, NaN, NaN, 1029.2523, 1029.2277, 1029.1914, 1029.1449, 1029.1038, 1029.0626, 1029.0184, 1028.9747, 1028.9247, 1028.868, 1028.8159, 1028.762, 1028.7091, 1028.6558, 1028.6082, 1028.5564, 1028.5045, 1028.4481, 1028.3984, 1028.3496, 1028.2949, 1028.2455, 1028.1951, 1028.1425, 1028.0823, 1028.0325, 1027.9786, 1027.9259, 1027.8735, 1027.8121, 1027.756, 1027.7056, 1027.6522, 1027.6012, 1027.5496, 1027.4857, 1027.4366, 1027.377, 1027.3083, 1027.2438, 1027.1757, 1027.1045, 1027.0359, 1026.9425, 1026.8176, 1026.6835, 1026.5013, 1026.3888, 1026.2148, 1026.0267, 1025.8761, 1025.7861, 1025.6667, 1025.463, 1025.323, 1025.252, 1025.1396, 1024.9802, 1024.7921, 1024.5806, 1024.4178, 1024.1868, 1024.112, 1024.0071, 1023.92676, 1023.86786, 1023.8365, 1023.81445, 1023.79065, 1023.7705, NaN, NaN, 1029.2366, 1029.2095, 1029.1685, 1029.1188, 1029.0703, 1029.0189, 1028.9677, 1028.919, 1028.8727, 1028.8229, 1028.7694, 1028.7188, 1028.6666, 1028.6133, 1028.5566, 1028.5044, 1028.4471, 1028.3912, 1028.333, 1028.2823, 1028.2312, 1028.1772, 1028.1243, 1028.0677, 1028.0105, 1027.9443, 1027.8853, 1027.8268, 1027.7698, 1027.718, 1027.6633, 1027.613, 1027.5563, 1027.499, 1027.4475, 1027.379, 1027.3126, 1027.2538, 1027.1836, 1027.1216, 1027.039, 1026.9302, 1026.819, 1026.7001, 1026.5939, 1026.4762, 1026.3682, 1026.2211, 1026.0472, 1025.9061, 1025.7252, 1025.5726, 1025.4865, 1025.32, 1025.192, 1025.0853, 1024.9716, 1024.728, 1024.4769, 1024.1917, 1024.1019, 1024.0369, 1023.9433, 1023.8641, 1023.8242, 1023.8027, 1023.77966, 1023.75555, 1023.7391, NaN, NaN, 1029.2499, 1029.2191, 1029.1819, 1029.1267, 1029.0757, 1029.019, 1028.9655, 1028.909, 1028.8549, 1028.7991, 1028.744, 1028.6901, 1028.6377, 1028.5885, 1028.5343, 1028.478, 1028.425, 1028.3741, 1028.3185, 1028.2584, 1028.2015, 1028.1456, 1028.0939, 1028.0386, 1027.9849, 1027.9293, 1027.8779, 1027.8243, 1027.7697, 1027.7136, 1027.6643, 1027.6079, 1027.5516, 1027.4833, 1027.4281, 1027.3699, 1027.314, 1027.2567, 1027.1787, 1027.0916, 1026.9974, 1026.9005, 1026.7804, 1026.6771, 1026.5759, 1026.4224, 1026.2965, 1026.1041, 1025.9797, 1025.822, 1025.702, 1025.5535, 1025.4695, 1025.3304, 1025.23, 1025.1255, 1025.0309, 1024.9448, 1024.8154, 1024.4845, 1024.186, 1024.0254, 1023.8771, 1023.8144, 1023.79016, 1023.7645, 1023.7302, 1023.70013, NaN, NaN, 1029.2483, 1029.2211, 1029.1855, 1029.1361, 1029.0931, 1029.0469, 1029.0002, 1028.9583, 1028.913, 1028.8668, 1028.8181, 1028.7684, 1028.7231, 1028.6737, 1028.625, 1028.5754, 1028.5309, 1028.4867, 1028.4359, 1028.388, 1028.3403, 1028.2941, 1028.2499, 1028.2028, 1028.1561, 1028.1094, 1028.0613, 1028.018, 1027.9641, 1027.9116, 1027.8506, 1027.7986, 1027.7472, 1027.6969, 1027.6477, 1027.5989, 1027.551, 1027.4913, 1027.4387, 1027.3824, 1027.3185, 1027.2529, 1027.1849, 1027.0947, 1027.0183, 1026.9216, 1026.8223, 1026.7062, 1026.6058, 1026.4786, 1026.3446, 1026.1803, 1026.0505, 1025.9155, 1025.733, 1025.5696, 1025.485, 1025.3616, 1025.2023, 1025.0592, 1024.9517, 1024.836, 1024.5692, 1024.2676, 1024.1327, 1024.0022, 1023.8846, 1023.82214, 1023.7852, 1023.74976, 1023.7163, 1023.6876, NaN, NaN, 1029.2576, 1029.2268, 1029.1893, 1029.1437, 1029.0996, 1029.0541, 1029.0093, 1028.9573, 1028.9027, 1028.8585, 1028.8092, 1028.7611, 1028.7162, 1028.6682, 1028.6172, 1028.5654, 1028.5173, 1028.468, 1028.414, 1028.3596, 1028.3112, 1028.2527, 1028.1884, 1028.1277, 1028.0682, 1028.0187, 1027.9653, 1027.9081, 1027.8567, 1027.8076, 1027.76, 1027.7059, 1027.6396, 1027.5765, 1027.5177, 1027.4703, 1027.4126, 1027.3423, 1027.2781, 1027.206, 1027.1288, 1027.0498, 1026.9691, 1026.8666, 1026.7451, 1026.5695, 1026.3832, 1026.2295, 1026.0857, 1025.9507, 1025.8193, 1025.6735, 1025.5444, 1025.4261, 1025.324, 1025.2137, 1025.0901, 1024.9949, 1024.8535, 1024.6276, 1024.5049, 1024.2601, 1024.0792, 1023.9061, 1023.8228, 1023.78406, 1023.758, 1023.7347, 1023.7137, 1023.70056, NaN, NaN, 1029.2594, 1029.2323, 1029.192, 1029.139, 1029.0891, 1029.0396, 1028.9802, 1028.9269, 1028.875, 1028.8219, 1028.7712, 1028.7213, 1028.6733, 1028.625, 1028.5734, 1028.5245, 1028.4792, 1028.4331, 1028.3828, 1028.3292, 1028.2761, 1028.2161, 1028.1641, 1028.104, 1028.0454, 1027.9889, 1027.9276, 1027.8694, 1027.8195, 1027.7576, 1027.7002, 1027.6499, 1027.595, 1027.5344, 1027.4746, 1027.4175, 1027.355, 1027.2919, 1027.2297, 1027.1562, 1027.0884, 1027.0103, 1026.9185, 1026.7947, 1026.6764, 1026.5157, 1026.3634, 1026.217, 1026.0381, 1025.9104, 1025.7885, 1025.6431, 1025.5269, 1025.3956, 1025.2426, 1025.1351, 1025.0238, 1024.8286, 1024.5878, 1024.3392, 1024.1427, 1024.0134, 1023.9055, 1023.7981, 1023.76935, 1023.7434, 1023.7114, 1023.6896, NaN, NaN, 1029.2609, 1029.2294, 1029.1932, 1029.1494, 1029.1066, 1029.0592, 1029.01, 1028.9615, 1028.9117, 1028.8602, 1028.809, 1028.7577, 1028.7069, 1028.6595, 1028.6079, 1028.5559, 1028.5071, 1028.4525, 1028.3984, 1028.3539, 1028.3013, 1028.2523, 1028.1984, 1028.1544, 1028.1073, 1028.056, 1028.0015, 1027.9504, 1027.8951, 1027.8457, 1027.7974, 1027.7423, 1027.684, 1027.6234, 1027.5724, 1027.5208, 1027.4664, 1027.4044, 1027.3341, 1027.2738, 1027.1995, 1027.1187, 1027.0258, 1026.926, 1026.8269, 1026.7542, 1026.6599, 1026.5297, 1026.373, 1026.2292, 1026.1025, 1025.9806, 1025.8463, 1025.6896, 1025.5771, 1025.4694, 1025.4016, 1025.3162, 1025.1854, 1025.12, 1025.0106, 1024.9099, 1024.759, 1024.5985, 1024.3531, 1024.0978, 1023.89777, 1023.84674, 1023.8112, 1023.79205, 1023.7694, 1023.75, NaN, NaN, 1029.2582, 1029.2303, 1029.1881, 1029.132, 1029.0808, 1029.0234, 1028.9648, 1028.9104, 1028.8602, 1028.8097, 1028.754, 1028.7054, 1028.6542, 1028.6042, 1028.5491, 1028.4962, 1028.4419, 1028.3817, 1028.3373, 1028.2844, 1028.2302, 1028.1803, 1028.1292, 1028.0763, 1028.0277, 1027.9763, 1027.9204, 1027.8683, 1027.8134, 1027.7559, 1027.7054, 1027.6505, 1027.5966, 1027.5437, 1027.4867, 1027.4348, 1027.3694, 1027.2946, 1027.2274, 1027.1738, 1027.1085, 1027.0171, 1026.9229, 1026.8198, 1026.7157, 1026.6292, 1026.5121, 1026.3926, 1026.2465, 1026.0677, 1025.9023, 1025.7701, 1025.6304, 1025.4811, 1025.3402, 1025.2478, 1025.1165, 1025.0474, 1024.9598, 1024.8579, 1024.7128, 1024.1627, 1023.9348, 1023.9072, 1023.87585, 1023.85425, 1023.8359, 1023.809, 1023.8006, NaN, NaN, 1029.2512, 1029.2251, 1029.1901, 1029.1498, 1029.108, 1029.0652, 1029.0178, 1028.9708, 1028.9204, 1028.8702, 1028.8223, 1028.7755, 1028.7264, 1028.6768, 1028.6295, 1028.5845, 1028.5314, 1028.4823, 1028.4297, 1028.3755, 1028.3179, 1028.2659, 1028.203, 1028.1556, 1028.1094, 1028.0603, 1028.0078, 1027.9537, 1027.9031, 1027.8553, 1027.8027, 1027.7559, 1027.7004, 1027.6449, 1027.5846, 1027.5306, 1027.4791, 1027.4135, 1027.3539, 1027.2955, 1027.2267, 1027.1422, 1027.0615, 1026.9983, 1026.9062, 1026.8011, 1026.6984, 1026.6135, 1026.5286, 1026.4221, 1026.2759, 1026.1682, 1025.984, 1025.841, 1025.7015, 1025.5703, 1025.4332, 1025.3082, 1025.1799, 1025.0814, 1024.9712, 1024.8704, 1024.6898, 1024.2511, 1023.99805, 1023.9696, 1023.94965, 1023.9259, 1023.90765, NaN, NaN, 1029.2767, 1029.2509, 1029.2144, 1029.1633, 1029.1163, 1029.0671, 1029.0178, 1028.9655, 1028.9133, 1028.8574, 1028.8064, 1028.7588, 1028.7007, 1028.6509, 1028.5979, 1028.5474, 1028.4962, 1028.4425, 1028.3898, 1028.3339, 1028.2784, 1028.2168, 1028.1571, 1028.1012, 1028.046, 1027.9905, 1027.9386, 1027.8848, 1027.8304, 1027.7812, 1027.7261, 1027.6681, 1027.6055, 1027.5509, 1027.4849, 1027.4276, 1027.3696, 1027.3086, 1027.2384, 1027.173, 1027.0936, 1027.0145, 1026.9473, 1026.8524, 1026.7494, 1026.6454, 1026.532, 1026.3921, 1026.2236, 1026.0715, 1025.8927, 1025.7848, 1025.6714, 1025.5376, 1025.3971, 1025.2418, 1025.0853, 1024.9738, 1024.8127, 1024.6682, 1024.4308, 1024.1886, 1024.0708, 1024.0396, 1024.0161, 1023.98376, NaN, NaN, 1029.27, 1029.2455, 1029.2147, 1029.175, 1029.1346, 1029.0848, 1029.0417, 1028.9946, 1028.9513, 1028.9038, 1028.8569, 1028.8143, 1028.7697, 1028.7263, 1028.6815, 1028.636, 1028.5916, 1028.5383, 1028.4902, 1028.4382, 1028.3839, 1028.329, 1028.2795, 1028.2306, 1028.1759, 1028.1238, 1028.0682, 1028.0135, 1027.9589, 1027.913, 1027.8612, 1027.8048, 1027.7498, 1027.6967, 1027.6456, 1027.5869, 1027.5275, 1027.4701, 1027.4175, 1027.3531, 1027.2855, 1027.2218, 1027.1516, 1027.07, 1026.9789, 1026.8923, 1026.7865, 1026.6853, 1026.5813, 1026.466, 1026.3369, 1026.1996, 1026.0256, 1025.8885, 1025.7643, 1025.6289, 1025.5149, 1025.4016, 1025.2964, 1025.1964, 1025.0972, 1024.994, 1024.9175, 1024.7782, 1024.6261, 1024.4192, 1024.0571, 1023.9557, 1023.9336, 1023.90936, 1023.8862, 1023.8661, NaN, NaN, 1029.2661, 1029.2393, 1029.2019, 1029.1526, 1029.0963, 1029.0444, 1028.9899, 1028.9341, 1028.8788, 1028.8254, 1028.769, 1028.7157, 1028.6583, 1028.6033, 1028.5514, 1028.4967, 1028.4424, 1028.3904, 1028.336, 1028.2864, 1028.2329, 1028.1802, 1028.1228, 1028.0742, 1028.0189, 1027.9609, 1027.898, 1027.839, 1027.7749, 1027.7094, 1027.6451, 1027.5933, 1027.525, 1027.461, 1027.3995, 1027.3353, 1027.2814, 1027.2186, 1027.1624, 1027.0883, 1027.0142, 1026.9441, 1026.8708, 1026.7703, 1026.6617, 1026.5428, 1026.3961, 1026.2178, 1026.0647, 1025.8911, 1025.7336, 1025.5734, 1025.433, 1025.3289, 1025.2144, 1025.1193, 1025.0054, 1024.9166, 1024.7626, 1024.6448, 1024.4014, 1024.0028, 1023.9495, 1023.86945, 1023.8296, 1023.8041, 1023.78973, NaN, NaN, 1029.2759, 1029.2437, 1029.2072, 1029.1578, 1029.1039, 1029.0498, 1029.0015, 1028.9498, 1028.8942, 1028.8346, 1028.7871, 1028.7401, 1028.6859, 1028.6311, 1028.5763, 1028.5195, 1028.4652, 1028.415, 1028.3591, 1028.3015, 1028.2526, 1028.1981, 1028.1426, 1028.0824, 1028.0248, 1027.9756, 1027.9192, 1027.8643, 1027.8075, 1027.7557, 1027.6912, 1027.6392, 1027.5901, 1027.5326, 1027.4813, 1027.425, 1027.3712, 1027.323, 1027.2639, 1027.1829, 1027.1118, 1027.0376, 1026.9569, 1026.8541, 1026.736, 1026.646, 1026.5366, 1026.4103, 1026.2323, 1025.9916, 1025.8379, 1025.7168, 1025.6389, 1025.5144, 1025.3964, 1025.2103, 1025.1052, 1025.0361, 1024.9594, 1024.7997, 1024.6229, 1024.245, 1024.0101, 1023.95416, 1023.91815, 1023.853, 1023.811, NaN, NaN, 1029.2571, 1029.23, 1029.1975, 1029.1469, 1029.1034, 1029.051, 1029.0033, 1028.9536, 1028.9005, 1028.8463, 1028.7911, 1028.7444, 1028.6924, 1028.6494, 1028.6062, 1028.5608, 1028.5125, 1028.4641, 1028.4244, 1028.3812, 1028.3334, 1028.2795, 1028.2292, 1028.1792, 1028.1322, 1028.0812, 1028.0295, 1027.9862, 1027.9375, 1027.888, 1027.8379, 1027.7906, 1027.7346, 1027.6779, 1027.6248, 1027.5762, 1027.5244, 1027.4628, 1027.3984, 1027.336, 1027.2919, 1027.2269, 1027.1633, 1027.0933, 1027.0194, 1026.9507, 1026.8749, 1026.7704, 1026.6569, 1026.5538, 1026.43, 1026.2653, 1026.0963, 1025.902, 1025.6853, 1025.5369, 1025.4246, 1025.3167, 1025.2258, 1025.1309, 1025.0461, 1024.9344, 1024.8086, 1024.629, 1024.2633, 1024.076, 1024.0447, 1024.0161, 1023.9579, 1023.89325, NaN, NaN, 1029.2526, 1029.227, 1029.1892, 1029.1392, 1029.0858, 1029.0338, 1028.9825, 1028.9357, 1028.8805, 1028.8341, 1028.7782, 1028.7355, 1028.69, 1028.6404, 1028.5858, 1028.5355, 1028.483, 1028.428, 1028.3768, 1028.3326, 1028.2815, 1028.2305, 1028.1772, 1028.1204, 1028.061, 1028.001, 1027.9418, 1027.8872, 1027.8326, 1027.7764, 1027.7299, 1027.6724, 1027.6178, 1027.5608, 1027.5006, 1027.4502, 1027.3949, 1027.332, 1027.271, 1027.2173, 1027.1648, 1027.109, 1027.0408, 1026.9705, 1026.8823, 1026.7963, 1026.6636, 1026.5823, 1026.4768, 1026.3328, 1026.183, 1026.0504, 1025.9448, 1025.8074, 1025.6586, 1025.4274, 1025.3226, 1025.1898, 1025.0806, 1024.8499, 1024.7238, 1024.3971, 1024.0339, 1023.98694, 1023.97076, 1023.94165, 1023.9255, NaN, NaN, 1029.2837, 1029.2587, 1029.2177, 1029.1683, 1029.1205, 1029.0685, 1029.0201, 1028.9717, 1028.925, 1028.8754, 1028.8167, 1028.7739, 1028.7242, 1028.6748, 1028.6324, 1028.5828, 1028.5364, 1028.4897, 1028.4382, 1028.3798, 1028.3253, 1028.2781, 1028.2234, 1028.1741, 1028.1232, 1028.0746, 1028.0208, 1027.9735, 1027.9238, 1027.8711, 1027.8198, 1027.7722, 1027.7222, 1027.6724, 1027.6224, 1027.5691, 1027.5117, 1027.4622, 1027.4143, 1027.363, 1027.3029, 1027.2307, 1027.1448, 1027.0812, 1027.0032, 1026.9231, 1026.8385, 1026.7632, 1026.649, 1026.5317, 1026.3646, 1026.2275, 1026.0741, 1025.9119, 1025.7516, 1025.5679, 1025.4564, 1025.3386, 1025.1846, 1024.9937, 1024.879, 1024.6931, 1024.5048, 1024.2733, 1024.0208, 1023.974, 1023.9525, 1023.93555, NaN, NaN, 1029.2606, 1029.2366, 1029.2021, 1029.1566, 1029.1116, 1029.0618, 1029.0079, 1028.9556, 1028.8978, 1028.841, 1028.7834, 1028.7349, 1028.6863, 1028.6313, 1028.5759, 1028.5242, 1028.4751, 1028.4249, 1028.3712, 1028.3232, 1028.272, 1028.226, 1028.1711, 1028.1077, 1028.0537, 1028.0107, 1027.957, 1027.8986, 1027.8458, 1027.8003, 1027.7526, 1027.7057, 1027.6478, 1027.5936, 1027.5404, 1027.4905, 1027.4392, 1027.3888, 1027.3281, 1027.2811, 1027.229, 1027.1682, 1027.1116, 1027.0524, 1026.9806, 1026.9036, 1026.8304, 1026.7357, 1026.6188, 1026.5402, 1026.4064, 1026.231, 1026.0867, 1025.9188, 1025.7836, 1025.6853, 1025.5227, 1025.3741, 1025.2417, 1025.0686, 1024.8987, 1024.7794, 1024.6187, 1024.5057, 1024.2468, 1024.0781, 1023.9518, 1023.8874, 1023.87274, NaN, NaN, 1029.2734, 1029.2313, 1029.1913, 1029.1481, 1029.1006, 1029.0426, 1028.9976, 1028.9534, 1028.9115, 1028.859, 1028.8196, 1028.7811, 1028.729, 1028.6752, 1028.6204, 1028.5651, 1028.516, 1028.4688, 1028.4194, 1028.3612, 1028.303, 1028.2501, 1028.2032, 1028.1506, 1028.0913, 1028.0353, 1027.9873, 1027.9346, 1027.8817, 1027.8254, 1027.7673, 1027.7092, 1027.6595, 1027.6077, 1027.5458, 1027.4968, 1027.4459, 1027.3931, 1027.3324, 1027.2812, 1027.2196, 1027.1599, 1027.1007, 1027.0319, 1026.9706, 1026.9043, 1026.8315, 1026.7238, 1026.6287, 1026.5482, 1026.4235, 1026.3514, 1026.225, 1026.1089, 1025.956, 1025.8102, 1025.6418, 1025.5214, 1025.4515, 1025.3951, 1025.34, 1025.2048, 1024.9407, 1024.8418, 1024.7274, 1024.6246, 1024.4812, 1024.096, 1023.9033, 1023.8855, NaN, NaN, 1029.2748, 1029.2422, 1029.1981, 1029.1431, 1029.0956, 1029.0514, 1029.0009, 1028.9552, 1028.9086, 1028.859, 1028.8114, 1028.771, 1028.7198, 1028.6626, 1028.607, 1028.5544, 1028.5073, 1028.4563, 1028.4149, 1028.3657, 1028.3127, 1028.2645, 1028.2076, 1028.1682, 1028.11, 1028.0544, 1028.0035, 1027.9581, 1027.8988, 1027.8511, 1027.8016, 1027.7534, 1027.7006, 1027.6365, 1027.5746, 1027.522, 1027.4608, 1027.4039, 1027.3474, 1027.2894, 1027.2333, 1027.1715, 1027.122, 1027.0596, 1027.0068, 1026.9546, 1026.8751, 1026.798, 1026.6554, 1026.5154, 1026.435, 1026.2827, 1026.135, 1025.9884, 1025.8516, 1025.7382, 1025.5785, 1025.4478, 1025.345, 1025.2578, 1025.1447, 1024.9896, 1024.8789, 1024.8151, 1024.7227, 1024.5632, 1024.0754, 1023.9331, 1023.92303, NaN, NaN, 1029.2175, 1029.1907, 1029.1554, 1029.0974, 1029.0435, 1028.9811, 1028.9272, 1028.8811, 1028.826, 1028.7719, 1028.715, 1028.6658, 1028.6099, 1028.556, 1028.5071, 1028.4607, 1028.4034, 1028.3401, 1028.2865, 1028.2268, 1028.1759, 1028.1183, 1028.069, 1028.0186, 1027.9636, 1027.9172, 1027.8606, 1027.7966, 1027.7325, 1027.6703, 1027.609, 1027.5645, 1027.5188, 1027.4609, 1027.3994, 1027.3518, 1027.3009, 1027.2498, 1027.1873, 1027.1277, 1027.0623, 1026.9873, 1026.9072, 1026.8285, 1026.7435, 1026.6888, 1026.617, 1026.5365, 1026.4485, 1026.308, 1026.1659, 1026.0258, 1025.9142, 1025.7662, 1025.5934, 1025.4761, 1025.338, 1025.149, 1024.9807, 1024.8403, 1024.7228, 1024.5427, 1024.172, 1024.0627, NaN, NaN, 1028.5465, 1028.5211, 1028.4893, 1028.4431, 1028.3854, 1028.3221, 1028.2609, 1028.1995, 1028.1521, 1028.096, 1028.0435, 1027.9993, 1027.9539, 1027.8999, 1027.8308, 1027.7726, 1027.7155, 1027.6642, 1027.6006, 1027.5314, 1027.4717, 1027.3986, 1027.3237, 1027.2611, 1027.2047, 1027.1488, 1027.0881, 1027.0231, 1026.939, 1026.8496, 1026.7616, 1026.6827, 1026.597, 1026.5262, 1026.4413, 1026.3801, 1026.3097, 1026.1803, 1026.075, 1025.9979, 1025.916, 1025.7156, 1025.4131, 1025.3232, 1025.2129, 1025.109, 1025.0414, 1024.9161, 1024.7416, 1024.5863, 1024.5085, NaN, NaN, 1028.2046, 1028.1708, 1028.1205, 1028.0476, 1027.9886, 1027.9288, 1027.8779, 1027.8318, 1027.7832, 1027.7289, 1027.6807, 1027.606, 1027.5321, 1027.4514, 1027.3922, 1027.3256, 1027.2428, 1027.1458, 1027.082, 1027.0243, 1026.9619, 1026.8838, 1026.8291, 1026.7402, 1026.6519, 1026.6019, 1026.5459, 1026.4238, 1026.2886, 1026.1364, 1026.0616, 1025.9724, 1025.8644, 1025.7969, 1025.5713, 1025.41, 1025.2291, 1025.0912, 1024.9974, 1024.8119, 1024.5905, 1024.4137, NaN, NaN, 1027.7557, 1027.7288, 1027.6624, 1027.5831, 1027.5265, 1027.4819, 1027.4423, 1027.3918, 1027.3278, 1027.2327, 1027.1755, 1027.1222, 1027.0586, 1027.0092, 1026.9479, 1026.87, 1026.8257, 1026.7533, 1026.6941, 1026.5845, 1026.4434, 1026.3026, 1026.2085, 1026.1454, 1026.068, 1025.9834, 1025.8619, 1025.6666, 1025.4498, 1025.2705, 1025.157, 1025.0364, 1024.8292, 1024.6599, 1024.4324, 1024.3323, NaN, NaN, 1027.312, 1027.2363, 1027.1759, 1027.099, 1027.0444, 1026.9912, 1026.9535, 1026.9111, 1026.8516, 1026.783, 1026.7019, 1026.6146, 1026.4812, 1026.2639, 1026.1583, 1026.0308, 1025.9231, 1025.852, 1025.7445, 1025.4949, 1025.2639, 1025.1453, 1024.9507, 1024.7672, 1024.6821, 1024.532, 1024.3439, NaN, NaN, 1027.2026, 1027.1609, 1027.1165, 1027.0498, 1026.9869, 1026.9359, 1026.8872, 1026.8298, 1026.7688, 1026.712, 1026.6265, 1026.5187, 1026.3755, 1026.1823, 1026.0331, 1025.9229, 1025.834, 1025.7296, 1025.5393, 1025.1677, 1025.0583, 1024.9211, 1024.7549, 1024.4003, 1024.3594, NaN, NaN, 1027.1509, 1027.1191, 1027.0815, 1027.0315, 1026.9683, 1026.9196, 1026.8745, 1026.8306, 1026.773, 1026.7109, 1026.6476, 1026.5817, 1026.4249, 1026.2312, 1026.0957, 1025.9473, 1025.8643, 1025.713, 1025.5427, 1025.2924, 1025.0237, 1024.762, 1024.5353, 1024.3649, NaN, NaN, 1027.1887, 1027.1423, 1027.1095, 1027.0691, 1027.0297, 1026.9819, 1026.9327, 1026.8816, 1026.8309, 1026.7798, 1026.718, 1026.6578, 1026.5342, 1026.4027, 1026.2184, 1026.132, 1026.004, 1025.8796, 1025.7051, 1025.5994, 1025.481, 1025.1683, 1024.8724, 1024.6423, 1024.4381, 1024.3806, NaN, NaN, 1027.1396, 1027.1091, 1027.0726, 1027.0072, 1026.9374, 1026.8867, 1026.8431, 1026.8004, 1026.7489, 1026.6768, 1026.5426, 1026.3661, 1026.2456, 1026.1598, 1026.0797, 1025.9152, 1025.6797, 1025.458, 1025.1614, 1024.8169, 1024.564, 1024.488, 1024.4402, NaN, NaN, 1027.1195, 1027.0847, 1027.0448, 1026.9752, 1026.9116, 1026.8494, 1026.7887, 1026.7299, 1026.621, 1026.4547, 1026.3331, 1026.2661, 1026.1852, 1026.1254, 1026.0642, 1025.9819, 1025.8721, 1025.7522, 1025.5518, 1025.3517, 1025.1212, 1024.8202, 1024.5555, 1024.4575, NaN, NaN, 1027.166, 1027.1221, 1027.0688, 1027.0195, 1026.9703, 1026.9225, 1026.8634, 1026.815, 1026.7643, 1026.7104, 1026.6544, 1026.6035, 1026.4559, 1026.2799, 1026.1711, 1026.1268, 1026.0718, 1026.0273, 1025.9464, 1025.8417, 1025.6943, 1025.4229, 1025.191, 1024.8937, 1024.7242, 1024.5267, 1024.4498, NaN, NaN, 1027.1804, 1027.1581, 1027.1313, 1027.092, 1027.0398, 1026.9594, 1026.9061, 1026.863, 1026.8114, 1026.7449, 1026.6918, 1026.6506, 1026.6017, 1026.5436, 1026.3911, 1026.2948, 1026.1888, 1026.1027, 1026.059, 1026.0034, 1025.9437, 1025.8701, 1025.7316, 1025.3833, 1024.9485, 1024.635, 1024.4836, NaN, NaN, 1027.0854, 1027.0521, 1027.0074, 1026.9457, 1026.8981, 1026.8474, 1026.7871, 1026.7184, 1026.6224, 1026.569, 1026.3829, 1026.2322, 1026.1539, 1026.0876, 1026.0365, 1025.9751, 1025.8916, 1025.7998, 1025.5452, 1025.145, 1024.667, 1024.5779, NaN, NaN, 1027.1063, 1027.0353, 1026.9812, 1026.9307, 1026.8832, 1026.839, 1026.792, 1026.7523, 1026.7029, 1026.6337, 1026.5844, 1026.512, 1026.4364, 1026.3141, 1026.215, 1026.1222, 1026.0688, 1025.9926, 1025.8916, 1025.7892, 1025.5614, 1025.367, 1025.2173, 1025.1166, 1024.7897, 1024.6517, 1024.6338, NaN, NaN, 1027.1006, 1027.0751, 1027.006, 1026.9377, 1026.8806, 1026.8242, 1026.7727, 1026.7034, 1026.6388, 1026.5032, 1026.3286, 1026.2086, 1026.149, 1026.0596, 1025.983, 1025.8988, 1025.7694, 1025.6111, 1025.287, 1025.083, 1024.8207, 1024.6493, NaN, NaN, 1027.2198, 1027.1556, 1026.9911, 1026.9166, 1026.8562, 1026.8104, 1026.7633, 1026.6965, 1026.6399, 1026.5785, 1026.4785, 1026.3461, 1026.277, 1026.2006, 1026.1035, 1026.0073, 1025.8999, 1025.7496, 1025.4916, 1025.2292, 1024.9799, 1024.7347, 1024.642, NaN, NaN, 1027.0161, 1026.9645, 1026.9199, 1026.8741, 1026.8217, 1026.7662, 1026.7169, 1026.6443, 1026.5891, 1026.4968, 1026.3785, 1026.2726, 1026.1735, 1026.0956, 1026.0371, 1025.9674, 1025.8577, 1025.7064, 1025.4603, 1025.1222, 1024.7958, 1024.6621, NaN, NaN, 1026.9381, 1026.901, 1026.8319, 1026.7759, 1026.7261, 1026.65, 1026.5862, 1026.5417, 1026.4878, 1026.3856, 1026.303, 1026.2079, 1026.1409, 1026.0634, 1025.9657, 1025.8501, 1025.7249, 1025.5875, 1025.3434, 1025.0215, 1024.7682, 1024.6536, NaN, NaN, 1026.9364, 1026.909, 1026.8367, 1026.7593, 1026.6825, 1026.6122, 1026.546, 1026.5012, 1026.4221, 1026.3221, 1026.2358, 1026.166, 1026.0435, 1025.958, 1025.8114, 1025.6296, 1025.3008, 1024.9515, 1024.7385, 1024.6661, 1024.6626, 1024.6692, NaN, NaN, 1026.973, 1026.8854, 1026.8059, 1026.716, 1026.6278, 1026.5564, 1026.5105, 1026.4595, 1026.4082, 1026.3269, 1026.2518, 1026.1348, 1026.0541, 1025.9674, 1025.8518, 1025.7568, 1025.5665, 1025.304, 1024.9308, 1024.6859, 1024.6428, NaN, NaN, 1026.8947, 1026.8695, 1026.8048, 1026.7142, 1026.6285, 1026.5333, 1026.4799, 1026.4318, 1026.3816, 1026.3124, 1026.1289, 1026.0211, 1025.9092, 1025.7665, 1025.5896, 1025.3749, 1025.1932, 1024.981, 1024.7073, 1024.646, 1024.6415, NaN, NaN, 1026.96, 1026.9081, 1026.8477, 1026.7603, 1026.676, 1026.5901, 1026.5099, 1026.4569, 1026.4062, 1026.3477, 1026.1971, 1026.0632, 1025.98, 1025.7822, 1025.5422, 1025.3536, 1025.2495, 1025.0151, 1024.826, 1024.633, NaN, NaN, 1026.9573, 1026.8958, 1026.8567, 1026.7644, 1026.6849, 1026.6194, 1026.5455, 1026.4796, 1026.4308, 1026.3899, 1026.3381, 1026.2231, 1026.1382, 1026.0514, 1025.9316, 1025.7095, 1025.4076, 1025.2173, 1024.9622, 1024.6981, 1024.6295, 1024.6259, NaN, NaN, 1026.8744, 1026.8079, 1026.7185, 1026.6254, 1026.5406, 1026.4912, 1026.4357, 1026.3615, 1026.2722, 1026.1924, 1026.0967, 1025.9938, 1025.9142, 1025.8292, 1025.6531, 1025.3862, 1025.2379, 1025.0352, 1024.8376, 1024.5762, NaN, NaN, 1026.9111, 1026.8767, 1026.8422, 1026.7977, 1026.7448, 1026.6322, 1026.5648, 1026.472, 1026.4093, 1026.3595, 1026.2755, 1026.156, 1026.0054, 1025.8844, 1025.7303, 1025.5985, 1025.4154, 1025.194, 1024.9323, 1024.7441, 1024.6205, NaN, NaN, 1026.8718, 1026.8374, 1026.7926, 1026.7291, 1026.6722, 1026.5962, 1026.5322, 1026.4852, 1026.4395, 1026.3691, 1026.3218, 1026.2734, 1026.182, 1026.0796, 1025.9138, 1025.6871, 1025.4473, 1025.0006, 1024.6185, NaN, NaN, 1026.871, 1026.8391, 1026.7916, 1026.7375, 1026.6687, 1026.6129, 1026.5431, 1026.4961, 1026.4524, 1026.3887, 1026.305, 1026.2166, 1026.1255, 1025.9552, 1025.8636, 1025.6561, 1025.2964, 1024.7827, 1024.5818, NaN, NaN, 1026.8203, 1026.7721, 1026.7357, 1026.6685, 1026.6046, 1026.5513, 1026.505, 1026.4629, 1026.4026, 1026.3276, 1026.2582, 1026.1969, 1026.1191, 1025.9744, 1025.8954, 1025.7789, 1025.5702, 1025.1512, 1024.7217, NaN, NaN, 1026.8584, 1026.8303, 1026.7904, 1026.7192, 1026.6423, 1026.582, 1026.5217, 1026.4755, 1026.4297, 1026.3809, 1026.3038, 1026.2361, 1026.1436, 1026.0374, 1025.8958, 1025.7375, 1025.5724, 1025.2599, 1024.9159, 1024.865, NaN, NaN, 1026.8376, 1026.7864, 1026.7365, 1026.6772, 1026.6156, 1026.5608, 1026.52, 1026.4773, 1026.4406, 1026.3984, 1026.3538, 1026.282, 1026.1904, 1026.0632, 1025.9309, 1025.8236, 1025.6704, 1025.5217, 1025.1229, NaN, NaN, 1026.8617, 1026.8423, 1026.7946, 1026.713, 1026.6447, 1026.5692, 1026.4829, 1026.4229, 1026.3673, 1026.3081, 1026.2393, 1026.1462, 1026.0027, 1025.8688, 1025.6746, 1025.4258, 1025.1788, 1025.1062, NaN, NaN, 1026.8276, 1026.7968, 1026.7533, 1026.679, 1026.6072, 1026.532, 1026.4669, 1026.42, 1026.3726, 1026.3031, 1026.2194, 1026.1426, 1026.0027, 1025.8838, 1025.7302, 1025.5922, 1025.3518, 1025.2262, NaN, NaN, 1026.7859, 1026.7415, 1026.672, 1026.6064, 1026.5138, 1026.4323, 1026.2809, 1026.1373, 1025.9459, 1025.8274, 1025.7523, 1025.7362, 1025.7107, 1025.6632, 1025.6096, 1025.5295, 1025.3749, 1025.2932, NaN, NaN, 1026.746, 1026.6781, 1026.6309, 1026.558, 1026.4807, 1026.4097, 1026.3114, 1026.1627, 1026.08, 1025.9656, 1025.8651, 1025.785, 1025.7341, 1025.6562, 1025.4958, 1025.3972, 1025.3679, NaN, NaN, 1026.6953, 1026.6525, 1026.6049, 1026.5444, 1026.491, 1026.4309, 1026.3628, 1026.2524, 1026.1449, 1026.065, 1025.9349, 1025.8658, 1025.8275, 1025.784, 1025.726, 1025.6697, 1025.6055, 1025.4369, 1025.3545, NaN, NaN, 1026.7029, 1026.6532, 1026.6018, 1026.54, 1026.4513, 1026.3523, 1026.2297, 1026.1276, 1026.019, 1025.9104, 1025.7968, 1025.7153, 1025.64, 1025.5325, 1025.3953, 1025.3193, NaN, NaN, 1026.6864, 1026.6504, 1026.6152, 1026.5603, 1026.5054, 1026.4537, 1026.3936, 1026.3162, 1026.2257, 1026.13, 1026.0428, 1025.9539, 1025.8019, 1025.6871, 1025.6053, 1025.5065, 1025.4209, 1025.3335, 1025.3097, NaN, NaN, 1026.7363, 1026.7128, 1026.6727, 1026.5793, 1026.4979, 1026.3914, 1026.266, 1026.186, 1026.101, 1026.0372, 1025.9116, 1025.7831, 1025.6967, 1025.6361, 1025.5804, 1025.5089, 1025.3418, 1025.3226, 1025.3173, NaN, NaN, 1026.7292, 1026.7039, 1026.6691, 1026.6061, 1026.5232, 1026.3787, 1026.2316, 1026.1154, 1026.0404, 1025.962, 1025.8131, 1025.7039, 1025.6465, 1025.5779, 1025.4353, 1025.3325, NaN, NaN, 1026.7249, 1026.7002, 1026.6716, 1026.6295, 1026.584, 1026.5034, 1026.412, 1026.292, 1026.1555, 1026.0442, 1025.956, 1025.8745, 1025.7695, 1025.6659, 1025.5591, 1025.4552, 1025.4182, 1025.4099, 1025.4114, NaN, NaN, 1026.7041, 1026.6783, 1026.6472, 1026.6117, 1026.5721, 1026.5187, 1026.4263, 1026.3195, 1026.2019, 1026.0927, 1025.9906, 1025.8125, 1025.7478, 1025.666, 1025.5437, 1025.4366, 1025.4208, 1025.4208, NaN, NaN, 1026.7006, 1026.6802, 1026.6525, 1026.6139, 1026.5726, 1026.5114, 1026.4506, 1026.3529, 1026.2826, 1026.199, 1026.0994, 1025.943, 1025.8251, 1025.7528, 1025.6707, 1025.5328, 1025.4021, NaN, NaN, 1026.6982, 1026.6764, 1026.6462, 1026.6016, 1026.5453, 1026.4543, 1026.3495, 1026.2472, 1026.1232, 1025.974, 1025.8519, 1025.7628, 1025.6577, 1025.5131, 1025.3815, 1025.3607, 1025.357, NaN, NaN, 1026.6956, 1026.6733, 1026.6411, 1026.5931, 1026.5459, 1026.4836, 1026.3976, 1026.2831, 1026.1538, 1025.98, 1025.8577, 1025.7323, 1025.6443, 1025.4427, 1025.3073, 1025.2914, 1025.2882, NaN, NaN, 1026.662, 1026.6384, 1026.6097, 1026.5696, 1026.5206, 1026.4536, 1026.3663, 1026.286, 1026.1809, 1026.0608, 1025.9467, 1025.8557, 1025.7181, 1025.6124, 1025.4673, 1025.2411, NaN, NaN, 1026.6642, 1026.639, 1026.6056, 1026.5555, 1026.5029, 1026.4233, 1026.3412, 1026.2495, 1026.1294, 1025.9993, 1025.9011, 1025.7083, 1025.5526, 1025.2344, 1025.1841, 1025.1758, NaN, NaN, 1026.6285, 1026.605, 1026.5702, 1026.5245, 1026.4688, 1026.405, 1026.3433, 1026.248, 1026.152, 1026.0591, 1025.946, 1025.7504, 1025.567, 1025.2833, 1025.1733, NaN, NaN, 1026.6012, 1026.5752, 1026.5404, 1026.4894, 1026.4232, 1026.358, 1026.2854, 1026.2021, 1026.08, 1025.9752, 1025.841, 1025.6202, 1025.3107, NaN, NaN, 1026.622, 1026.5995, 1026.5691, 1026.5249, 1026.4783, 1026.4358, 1026.357, 1026.2896, 1026.188, 1026.1162, 1025.9899, 1025.8699, 1025.7341, 1025.554, 1025.3845, 1025.3187, 1025.314, NaN, NaN, 1026.5939, 1026.5685, 1026.5382, 1026.4973, 1026.4574, 1026.4031, 1026.3273, 1026.2825, 1026.2384, 1026.1735, 1026.0675, 1025.9843, 1025.8395, 1025.7598, 1025.5208, 1025.3704, 1025.3514, NaN, NaN, 1026.5784, 1026.5574, 1026.5251, 1026.4858, 1026.4481, 1026.4083, 1026.3589, 1026.2623, 1026.1741, 1026.073, 1025.9257, 1025.7997, 1025.6536, 1025.3512, NaN, NaN, 1026.5717, 1026.5458, 1026.5131, 1026.4705, 1026.4291, 1026.3572, 1026.2544, 1026.1327, 1026.0201, 1025.8661, 1025.7465, 1025.6221, 1025.336, 1025.2793, 1025.2711, NaN, NaN, 1026.5665, 1026.543, 1026.5151, 1026.4685, 1026.4128, 1026.3274, 1026.257, 1026.1631, 1026.0728, 1025.9365, 1025.7919, 1025.6886, 1025.5469, 1025.3619, 1025.3064, 1025.3096, NaN, NaN, 1026.5481, 1026.5248, 1026.4949, 1026.4557, 1026.4136, 1026.3602, 1026.2727, 1026.1705, 1026.0613, 1025.9763, 1025.7949, 1025.6459, 1025.5018, 1025.3297, NaN, NaN, 1026.5488, 1026.5262, 1026.4973, 1026.4584, 1026.4207, 1026.381, 1026.3097, 1026.2386, 1026.1427, 1025.997, 1025.8126, 1025.6055, 1025.4818, 1025.3555, 1025.2809, 1025.2814, NaN, NaN, 1026.5298, 1026.5032, 1026.4703, 1026.4296, 1026.384, 1026.3055, 1026.2216, 1026.0977, 1025.9648, 1025.7966, 1025.6179, 1025.4309, 1025.3392, 1025.3053, NaN, NaN, 1026.532, 1026.5084, 1026.4774, 1026.4346, 1026.3898, 1026.3428, 1026.2687, 1026.1302, 1026.026, 1025.8794, 1025.7407, 1025.5741, 1025.4248, NaN, NaN, 1026.5253, 1026.5046, 1026.4745, 1026.4357, 1026.3994, 1026.3618, 1026.3218, 1026.2657, 1026.1426, 1026.0394, 1025.9429, 1025.8038, 1025.644, 1025.5175, 1025.3866, 1025.3533, 1025.3492, NaN, NaN, 1026.493, 1026.4707, 1026.4396, 1026.395, 1026.3506, 1026.2972, 1026.1676, 1026.0408, 1025.9182, 1025.7311, 1025.5872, 1025.4232, 1025.3525, 1025.3362, 1025.3315, NaN, NaN, 1026.473, 1026.4467, 1026.4147, 1026.3756, 1026.3411, 1026.2865, 1026.1411, 1026.0316, 1025.8956, 1025.691, 1025.5552, 1025.4341, 1025.3507, NaN, NaN, 1026.4689, 1026.4443, 1026.4117, 1026.3643, 1026.3169, 1026.2267, 1026.0753, 1025.9596, 1025.7698, 1025.5927, 1025.4375, 1025.3784, 1025.3549, 1025.3433, NaN, NaN, 1026.4625, 1026.4391, 1026.4066, 1026.3712, 1026.3307, 1026.2428, 1026.1024, 1025.9714, 1025.8108, 1025.694, 1025.5493, 1025.4326, 1025.3761, 1025.3384, 1025.325, NaN, NaN, 1026.4414, 1026.418, 1026.3827, 1026.3389, 1026.2603, 1026.1002, 1025.9907, 1025.8381, 1025.7117, 1025.6127, 1025.4634, 1025.3668, 1025.3003, NaN, NaN, 1026.4136, 1026.3896, 1026.3593, 1026.3182, 1026.256, 1026.1188, 1025.9843, 1025.8495, 1025.6896, 1025.5863, 1025.4401, 1025.3602, 1025.3317, NaN, NaN, 1026.4335, 1026.4128, 1026.3855, 1026.3457, 1026.3027, 1026.2349, 1026.0872, 1025.975, 1025.8198, 1025.6818, 1025.5687, 1025.4576, 1025.4032, 1025.3562, 1025.3333, NaN, NaN, 1026.4186, 1026.3969, 1026.3644, 1026.3136, 1026.2202, 1026.0714, 1025.9305, 1025.734, 1025.6354, 1025.4937, 1025.392, NaN, NaN, 1026.408, 1026.3835, 1026.3534, 1026.3041, 1026.2112, 1026.0757, 1025.9207, 1025.751, 1025.6654, 1025.5343, 1025.4205, 1025.3167, 1025.3082, NaN, NaN, 1026.3989, 1026.3757, 1026.3467, 1026.2562, 1026.105, 1025.9365, 1025.787, 1025.716, 1025.6534, 1025.5356, 1025.4167, 1025.3033, 1025.2781, NaN, NaN, 1026.4036, 1026.3832, 1026.3516, 1026.3157, 1026.204, 1026.0936, 1025.9863, 1025.8394, 1025.7579, 1025.7075, 1025.5953, 1025.5197, 1025.4375, 1025.3123, 1025.2521, NaN, NaN, 1026.3856, 1026.3601, 1026.3242, 1026.1685, 1026.0308, 1025.9103, 1025.7709, 1025.7072, 1025.5963, 1025.4766, 1025.3315, 1025.2867, 1025.281, 1025.2799, NaN, NaN, 1026.4144, 1026.3984, 1026.3727, 1026.2911, 1026.1901, 1026.1185, 1026.0359, 1025.9227, 1025.8307, 1025.7291, 1025.6549, 1025.5563, 1025.361, 1025.303, 1025.3032, NaN, NaN, 1026.4296, 1026.4086, 1026.3795, 1026.343, 1026.3041, 1026.2357, 1026.1382, 1026.0839, 1025.9966, 1025.7618, 1025.6586, 1025.5127, 1025.2861, NaN, NaN, 1026.4572, 1026.4323, 1026.3953, 1026.3513, 1026.314, 1026.2692, 1026.2257, 1026.1508, 1026.0103, 1025.7461, 1025.6428, 1025.441, 1025.2512, 1025.241, NaN, NaN, 1026.4996, 1026.473, 1026.4369, 1026.3798, 1026.3252, 1026.2756, 1026.2305, 1026.1067, 1025.9342, 1025.6953, 1025.5779, 1025.3164, 1025.2383, 1025.2352, NaN, NaN, 1026.5464, 1026.5203, 1026.4893, 1026.4521, 1026.4171, 1026.3657, 1026.254, 1026.1642, 1026.0729, 1025.9543, 1025.7728, 1025.6539, 1025.4337, 1025.2358, NaN, NaN, 1026.5657, 1026.5421, 1026.5127, 1026.4729, 1026.4347, 1026.3573, 1026.1736, 1025.9912, 1025.8907, 1025.8336, 1025.771, 1025.7017, 1025.6238, 1025.3771, 1025.2599, 1025.2579, NaN, NaN, 1026.5964, 1026.5747, 1026.5464, 1026.5099, 1026.4675, 1026.4213, 1026.3572, 1026.239, 1026.108, 1025.8118, 1025.7246, 1025.6647, 1025.5822, 1025.4056, 1025.312, 1025.308, NaN, NaN, 1026.6278, 1026.607, 1026.5757, 1026.5398, 1026.5, 1026.4517, 1026.407, 1026.3335, 1026.1807, 1026.0288, 1025.817, 1025.6945, 1025.6384, 1025.5673, 1025.4004, 1025.3612, NaN, NaN, 1026.6561, 1026.636, 1026.6083, 1026.5634, 1026.519, 1026.4768, 1026.4363, 1026.3801, 1026.2279, 1026.092, 1025.8625, 1025.7592, 1025.6776, 1025.5934, 1025.4625, 1025.3903, 1025.383, NaN, NaN, 1026.6809, 1026.6592, 1026.6278, 1026.5862, 1026.5325, 1026.4285, 1026.3129, 1026.1692, 1026.0321, 1025.9099, 1025.8179, 1025.724, 1025.6241, 1025.5165, 1025.452, 1025.4338, 1025.4316, NaN, NaN, 1026.6884, 1026.6598, 1026.628, 1026.5902, 1026.5461, 1026.5006, 1026.4366, 1026.3683, 1026.232, 1026.0878, 1025.9417, 1025.8647, 1025.7709, 1025.6497, 1025.5267, 1025.464, NaN, NaN, 1026.698, 1026.6747, 1026.648, 1026.604, 1026.564, 1026.5217, 1026.4604, 1026.4095, 1026.3379, 1026.2544, 1026.0468, 1025.834, 1025.7264, 1025.5773, 1025.481, 1025.4384, 1025.427, 1025.428, NaN, NaN, 1026.7113, 1026.6888, 1026.6605, 1026.6215, 1026.5834, 1026.5391, 1026.4786, 1026.4048, 1026.3185, 1026.2457, 1026.1907, 1026.0742, 1025.8864, 1025.7324, 1025.546, 1025.4185, 1025.3875, 1025.378, NaN, NaN, 1026.7268, 1026.7035, 1026.675, 1026.6266, 1026.5801, 1026.5227, 1026.4657, 1026.3904, 1026.2551, 1026.1571, 1026.0504, 1025.9427, 1025.8276, 1025.6978, 1025.4617, 1025.3605, NaN, NaN, 1026.8741, 1026.8059, 1026.7578, 1026.7051, 1026.6619, 1026.6112, 1026.5579, 1026.4761, 1026.3536, 1026.2126, 1026.0648, 1025.9689, 1025.8616, 1025.7651, 1025.5951, 1025.3909, 1025.3025, 1025.2844, 1025.2808, NaN, NaN, 1026.8326, 1026.7714, 1026.7258, 1026.6691, 1026.6039, 1026.5531, 1026.4744, 1026.339, 1026.1606, 1026.0487, 1025.9069, 1025.8054, 1025.7037, 1025.6385, 1025.4952, 1025.324, 1025.1569, 1025.1403, 1025.1375, NaN, NaN, 1026.9248, 1026.866, 1026.8, 1026.7385, 1026.6614, 1026.612, 1026.5565, 1026.5028, 1026.4547, 1026.3916, 1026.3104, 1026.2579, 1026.1597, 1025.9669, 1025.7753, 1025.6317, 1025.3813, 1025.2211, 1025.0831, 1025.052, NaN, NaN, 1027.008, 1026.9775, 1026.9374, 1026.853, 1026.732, 1026.6632, 1026.5999, 1026.5294, 1026.4656, 1026.4104, 1026.3292, 1026.2627, 1026.1584, 1026.0311, 1025.8645, 1025.6967, 1025.4613, 1025.1731, 1024.9849, 1024.9614, 1024.9575, NaN, NaN, 1026.9769, 1026.9113, 1026.8696, 1026.7551, 1026.6886, 1026.6381, 1026.5891, 1026.519, 1026.4485, 1026.349, 1026.2728, 1026.1708, 1026.025, 1025.86, 1025.6865, 1025.4186, 1025.061, 1024.8922, 1024.8523, NaN, NaN, 1027.0309, 1026.9802, 1026.9181, 1026.8488, 1026.7732, 1026.7235, 1026.6819, 1026.6141, 1026.5406, 1026.4634, 1026.3942, 1026.3286, 1026.2686, 1026.1506, 1025.9761, 1025.8942, 1025.7749, 1025.6326, 1025.3546, 1024.985, 1024.8221, 1024.7968, 1024.7876, 1024.7891, NaN, NaN, 1027.0431, 1027.002, 1026.943, 1026.8608, 1026.8127, 1026.7477, 1026.651, 1026.603, 1026.5469, 1026.5016, 1026.4299, 1026.3292, 1026.2296, 1026.1147, 1025.9972, 1025.8909, 1025.8195, 1025.6357, 1025.4269, 1025.0891, 1024.823, 1024.7703, 1024.7456, NaN, NaN, 1027.0884, 1027.0437, 1026.9991, 1026.9275, 1026.8544, 1026.8022, 1026.7455, 1026.682, 1026.6084, 1026.5238, 1026.4774, 1026.4066, 1026.3184, 1026.2129, 1026.1406, 1026.0497, 1025.9185, 1025.707, 1025.4552, 1025.1359, 1024.8441, 1024.7441, 1024.7139, 1024.704, NaN, NaN, 1027.1276, 1027.0975, 1027.0312, 1026.9746, 1026.9086, 1026.848, 1026.7878, 1026.7272, 1026.6439, 1026.5729, 1026.496, 1026.4435, 1026.366, 1026.2736, 1026.209, 1026.1, 1025.8256, 1025.6465, 1025.5043, 1025.2812, 1024.9176, 1024.7489, 1024.7053, 1024.6663, NaN, NaN, 1027.2219, 1027.1824, 1027.0955, 1027.0271, 1026.9473, 1026.8945, 1026.8346, 1026.7667, 1026.7085, 1026.6399, 1026.5701, 1026.5151, 1026.4285, 1026.2925, 1026.2211, 1026.0963, 1025.8881, 1025.7308, 1025.5513, 1025.4072, 1025.1462, 1024.846, 1024.7411, 1024.6251, 1024.4944, 1024.4783, NaN, NaN, 1027.2987, 1027.2474, 1027.153, 1027.0901, 1027.0115, 1026.9403, 1026.8857, 1026.8315, 1026.7377, 1026.6042, 1026.531, 1026.4646, 1026.3861, 1026.3234, 1026.263, 1026.1945, 1026.0856, 1025.8522, 1025.6774, 1025.5055, 1025.3015, 1024.9717, 1024.7526, 1024.6633, 1024.3651, 1024.1068, NaN, NaN, 1027.2404, 1027.1774, 1027.1256, 1027.0475, 1026.9753, 1026.9122, 1026.834, 1026.7734, 1026.7207, 1026.6091, 1026.539, 1026.4601, 1026.3832, 1026.3113, 1026.1721, 1025.9978, 1025.8379, 1025.5636, 1025.3961, 1025.1807, 1024.9296, 1024.8726, 1024.7346, 1024.3484, 1024.0575, NaN, NaN, 1027.2871, 1027.2017, 1027.1566, 1027.1017, 1027.0397, 1026.9731, 1026.9081, 1026.8474, 1026.7928, 1026.7356, 1026.6884, 1026.6056, 1026.5005, 1026.3901, 1026.3271, 1026.2183, 1026.0553, 1025.8799, 1025.6924, 1025.5333, 1025.3446, 1025.0927, 1025.0013, 1024.7246, 1024.3885, 1024.1095, 1024.0632, NaN, NaN, 1027.4058, 1027.3707, 1027.3281, 1027.2743, 1027.2183, 1027.1495, 1027.0598, 1026.998, 1026.9369, 1026.8832, 1026.8397, 1026.7529, 1026.6938, 1026.6383, 1026.5237, 1026.4417, 1026.339, 1026.2262, 1026.0448, 1025.8387, 1025.607, 1025.4186, 1025.2603, 1025.1531, 1025.019, 1024.6897, 1024.3053, 1024.2032, 1024.0815, NaN, NaN, 1027.7745, 1027.7406, 1027.6808, 1027.61, 1027.5488, 1027.4797, 1027.4164, 1027.3704, 1027.329, 1027.2665, 1027.1588, 1027.0737, 1026.9879, 1026.9066, 1026.8334, 1026.7699, 1026.7219, 1026.67, 1026.5876, 1026.4615, 1026.3019, 1026.1445, 1026.0033, 1025.8623, 1025.727, 1025.5913, 1025.4606, 1025.2626, 1025.149, 1024.9607, 1024.6655, 1024.2825, 1024.1719, 1024.1519, NaN, NaN, 1028.2354, 1028.2115, 1028.1666, 1028.1089, 1028.0743, 1028.029, 1027.9728, 1027.9077, 1027.8523, 1027.813, 1027.7765, 1027.7175, 1027.6577, 1027.5988, 1027.547, 1027.4995, 1027.4269, 1027.3658, 1027.2786, 1027.1577, 1027.0879, 1027.0289, 1026.978, 1026.9044, 1026.8254, 1026.7645, 1026.6865, 1026.5947, 1026.493, 1026.374, 1026.245, 1026.0961, 1025.9446, 1025.7687, 1025.5895, 1025.3466, 1025.1327, 1024.9806, 1024.8339, 1024.6384, 1024.3522, 1024.2069, 1024.1707, 1024.1519, NaN, NaN, 1028.5829, 1028.5261, 1028.4961, 1028.4609, 1028.4263, 1028.3865, 1028.3457, 1028.2919, 1028.2456, 1028.2003, 1028.1484, 1028.0948, 1028.0415, 1027.9736, 1027.9208, 1027.8667, 1027.8177, 1027.7561, 1027.7039, 1027.658, 1027.6008, 1027.5421, 1027.4978, 1027.4506, 1027.3762, 1027.3066, 1027.2452, 1027.1959, 1027.1414, 1027.0809, 1027.0249, 1026.949, 1026.8574, 1026.781, 1026.6887, 1026.6113, 1026.5139, 1026.3956, 1026.2993, 1026.1969, 1026.0619, 1025.9364, 1025.7161, 1025.481, 1025.3348, 1025.1809, 1024.9767, 1024.7996, 1024.5258, 1024.269, 1024.1753, 1024.1466, 1024.1344, NaN, NaN, 1029.0885, 1029.0532, 1029.0184, 1028.9734, 1028.9338, 1028.8799, 1028.8267, 1028.7802, 1028.7247, 1028.6743, 1028.6265, 1028.5862, 1028.5477, 1028.5043, 1028.4564, 1028.4122, 1028.3594, 1028.3058, 1028.2582, 1028.2118, 1028.1594, 1028.1096, 1028.0604, 1028.0076, 1027.9602, 1027.9125, 1027.8673, 1027.821, 1027.7793, 1027.7296, 1027.6837, 1027.6315, 1027.5847, 1027.5375, 1027.4856, 1027.4388, 1027.3909, 1027.3408, 1027.287, 1027.2207, 1027.1702, 1027.1001, 1027.0421, 1026.9945, 1026.9458, 1026.8767, 1026.7921, 1026.724, 1026.6184, 1026.505, 1026.4025, 1026.2977, 1026.2351, 1026.1064, 1025.9939, 1025.7574, 1025.5991, 1025.4834, 1025.3787, 1025.2745, 1025.1753, 1025.0636, 1024.9133, 1024.7712, 1024.433, 1024.1892, 1024.1598, 1024.144, NaN, NaN, 1029.2721, 1029.2417, 1029.2119, 1029.1682, 1029.1101, 1029.0486, 1028.9987, 1028.9457, 1028.8994, 1028.8529, 1028.8007, 1028.7513, 1028.7037, 1028.6576, 1028.609, 1028.5613, 1028.5096, 1028.4591, 1028.4028, 1028.3541, 1028.3047, 1028.2548, 1028.2039, 1028.1532, 1028.1033, 1028.0513, 1027.9907, 1027.9264, 1027.8622, 1027.8105, 1027.7638, 1027.7118, 1027.6587, 1027.6014, 1027.5496, 1027.4949, 1027.4358, 1027.3788, 1027.3319, 1027.2676, 1027.1971, 1027.1296, 1027.0651, 1027.0074, 1026.9263, 1026.8441, 1026.7374, 1026.614, 1026.5236, 1026.4215, 1026.3362, 1026.1907, 1026.0444, 1025.9274, 1025.7732, 1025.6809, 1025.5267, 1025.3511, 1025.2302, 1025.1211, 1025.0393, 1024.933, 1024.6989, 1024.652, 1024.5614, 1024.3861, 1024.2694, 1024.2233, NaN, NaN, 1029.2665, 1029.2417, 1029.2059, 1029.1567, 1029.1093, 1029.0645, 1029.0154, 1028.9628, 1028.9144, 1028.8645, 1028.8181, 1028.7661, 1028.7214, 1028.6721, 1028.6207, 1028.5662, 1028.5156, 1028.4642, 1028.4192, 1028.3682, 1028.3243, 1028.2742, 1028.2213, 1028.1697, 1028.1145, 1028.0625, 1028.0079, 1027.9502, 1027.893, 1027.8425, 1027.7944, 1027.7415, 1027.6777, 1027.619, 1027.5704, 1027.5145, 1027.4598, 1027.3945, 1027.3445, 1027.286, 1027.2335, 1027.167, 1027.1107, 1027.0385, 1026.9803, 1026.8918, 1026.7924, 1026.7072, 1026.6277, 1026.5486, 1026.4474, 1026.3013, 1026.1029, 1025.9797, 1025.8741, 1025.6509, 1025.4752, 1025.403, 1025.2574, 1025.1012, 1024.8956, 1024.7764, 1024.6351, 1024.5227, 1024.408, 1024.3682, 1024.343, NaN, NaN, 1029.2781, 1029.2528, 1029.2213, 1029.1797, 1029.1301, 1029.0769, 1029.0282, 1028.9822, 1028.9344, 1028.8867, 1028.8379, 1028.7844, 1028.7253, 1028.6743, 1028.6257, 1028.5792, 1028.5276, 1028.4791, 1028.4312, 1028.3784, 1028.3279, 1028.2734, 1028.2142, 1028.1555, 1028.0974, 1028.043, 1027.9899, 1027.9276, 1027.8711, 1027.826, 1027.7749, 1027.7264, 1027.6859, 1027.6334, 1027.5713, 1027.5022, 1027.4543, 1027.4037, 1027.3458, 1027.2975, 1027.2532, 1027.2006, 1027.1237, 1027.0638, 1026.9832, 1026.9113, 1026.8358, 1026.7582, 1026.6956, 1026.6179, 1026.5089, 1026.3741, 1026.2284, 1026.0856, 1025.9904, 1025.8057, 1025.5879, 1025.4547, 1025.2714, 1025.0994, 1024.9485, 1024.8372, 1024.7041, 1024.6425, 1024.5443, 1024.3556, 1024.2991, NaN, NaN, 1029.2797, 1029.2504, 1029.2094, 1029.1671, 1029.1309, 1029.0853, 1029.0377, 1028.9885, 1028.9476, 1028.9015, 1028.8533, 1028.803, 1028.7502, 1028.7052, 1028.6534, 1028.6068, 1028.5591, 1028.5111, 1028.4612, 1028.4034, 1028.349, 1028.2928, 1028.24, 1028.1884, 1028.1355, 1028.0885, 1028.0353, 1027.9869, 1027.9384, 1027.8815, 1027.8279, 1027.7755, 1027.724, 1027.6654, 1027.6099, 1027.5565, 1027.5034, 1027.4457, 1027.39, 1027.3412, 1027.2838, 1027.2206, 1027.1736, 1027.1099, 1027.029, 1026.9553, 1026.8479, 1026.7664, 1026.6891, 1026.6111, 1026.527, 1026.4233, 1026.2549, 1026.1562, 1026.101, 1025.9536, 1025.8293, 1025.7634, 1025.6211, 1025.436, 1025.2084, 1025.0299, 1024.904, 1024.733, 1024.6274, 1024.59, 1024.5536, 1024.5149, 1024.4916, NaN, NaN, 1029.2577, 1029.2307, 1029.1953, 1029.1523, 1029.0994, 1029.0408, 1028.9838, 1028.9327, 1028.8816, 1028.8345, 1028.7811, 1028.7299, 1028.6787, 1028.6244, 1028.5636, 1028.5078, 1028.4541, 1028.4003, 1028.3417, 1028.291, 1028.243, 1028.1927, 1028.1428, 1028.0964, 1028.0497, 1028.0021, 1027.954, 1027.9065, 1027.8524, 1027.7909, 1027.7205, 1027.6709, 1027.614, 1027.5647, 1027.5055, 1027.4576, 1027.4065, 1027.3575, 1027.3068, 1027.2507, 1027.1915, 1027.1292, 1027.0483, 1026.9692, 1026.9089, 1026.8553, 1026.7751, 1026.6667, 1026.5886, 1026.542, 1026.4207, 1026.3112, 1026.1785, 1026.03, 1025.8762, 1025.7544, 1025.6675, 1025.4882, 1025.3553, 1025.1929, 1025.076, 1024.979, 1024.85, 1024.6776, 1024.5985, 1024.5554, 1024.4055, NaN, NaN, 1029.2649, 1029.2352, 1029.2029, 1029.1555, 1029.1049, 1029.0654, 1029.0166, 1028.9741, 1028.9247, 1028.8801, 1028.8334, 1028.7877, 1028.7397, 1028.6843, 1028.6338, 1028.5857, 1028.5353, 1028.4808, 1028.4291, 1028.383, 1028.3398, 1028.2859, 1028.2343, 1028.18, 1028.1211, 1028.0747, 1028.0284, 1027.977, 1027.9146, 1027.864, 1027.8079, 1027.7535, 1027.7007, 1027.6466, 1027.6014, 1027.559, 1027.5055, 1027.443, 1027.396, 1027.3451, 1027.29, 1027.2474, 1027.1941, 1027.143, 1027.0717, 1026.9983, 1026.9404, 1026.857, 1026.7822, 1026.6924, 1026.619, 1026.5304, 1026.4293, 1026.3107, 1026.1392, 1026.0038, 1025.8596, 1025.7736, 1025.692, 1025.5942, 1025.4551, 1025.3076, 1025.17, 1025.0087, 1024.9119, 1024.7823, 1024.655, 1024.5427, 1024.357, 1024.3008, NaN, NaN, 1029.2886, 1029.2621, 1029.2266, 1029.1718, 1029.1167, 1029.0597, 1029.0038, 1028.9514, 1028.8944, 1028.8336, 1028.7771, 1028.7279, 1028.6718, 1028.6134, 1028.556, 1028.5034, 1028.4479, 1028.3994, 1028.348, 1028.3021, 1028.2598, 1028.2053, 1028.1516, 1028.1006, 1028.0396, 1027.9872, 1027.9238, 1027.8594, 1027.8143, 1027.7646, 1027.7114, 1027.6672, 1027.6223, 1027.5736, 1027.5206, 1027.471, 1027.4093, 1027.357, 1027.3024, 1027.2372, 1027.1614, 1027.0854, 1027.0044, 1026.9343, 1026.8679, 1026.7612, 1026.6735, 1026.5779, 1026.4763, 1026.3324, 1026.1571, 1026.0001, 1025.8296, 1025.7423, 1025.6525, 1025.4827, 1025.3425, 1025.2277, 1025.0337, 1024.8811, 1024.7305, 1024.5087, 1024.2684, 1024.0911, 1024.0608, NaN, NaN, 1029.2833, 1029.2562, 1029.2145, 1029.1614, 1029.1105, 1029.061, 1029.0162, 1028.9716, 1028.9264, 1028.8823, 1028.8318, 1028.7725, 1028.7223, 1028.6658, 1028.6144, 1028.5702, 1028.5182, 1028.4711, 1028.4207, 1028.376, 1028.3336, 1028.2896, 1028.2413, 1028.1853, 1028.127, 1028.0741, 1028.0181, 1027.9604, 1027.9113, 1027.8536, 1027.8022, 1027.7454, 1027.6978, 1027.6484, 1027.5938, 1027.5405, 1027.4817, 1027.4202, 1027.3641, 1027.3098, 1027.26, 1027.2032, 1027.14, 1027.071, 1027.003, 1026.863, 1026.767, 1026.695, 1026.5978, 1026.477, 1026.3359, 1026.2224, 1026.0819, 1025.9825, 1025.8821, 1025.778, 1025.5792, 1025.4275, 1025.229, 1025.0417, 1024.8635, 1024.6412, 1024.3867, 1024.2198, 1024.1226, 1024.0751, 1024.0479, NaN, NaN, 1029.2802, 1029.2549, 1029.2266, 1029.1787, 1029.1293, 1029.0815, 1029.0336, 1028.9867, 1028.9397, 1028.8903, 1028.8342, 1028.78, 1028.7286, 1028.6785, 1028.6249, 1028.5713, 1028.5242, 1028.4749, 1028.4198, 1028.3723, 1028.3259, 1028.275, 1028.223, 1028.1649, 1028.1068, 1028.0509, 1027.9938, 1027.9423, 1027.888, 1027.8383, 1027.7927, 1027.7454, 1027.6929, 1027.6489, 1027.6011, 1027.5491, 1027.4886, 1027.4456, 1027.3958, 1027.339, 1027.2755, 1027.2198, 1027.1584, 1027.0939, 1027.0134, 1026.9438, 1026.8483, 1026.7983, 1026.725, 1026.6349, 1026.5333, 1026.3998, 1026.2461, 1026.086, 1025.9264, 1025.858, 1025.7211, 1025.5933, 1025.4515, 1025.3279, 1025.2112, 1025.0991, 1025.015, 1024.8868, 1024.7808, 1024.5157, 1024.1332, 1024.0874, 1024.0686, 1024.0518, NaN, NaN, 1029.2717, 1029.2445, 1029.209, 1029.1658, 1029.1233, 1029.0626, 1029.0142, 1028.9606, 1028.9135, 1028.8607, 1028.8127, 1028.7592, 1028.704, 1028.6562, 1028.6139, 1028.5675, 1028.5173, 1028.4666, 1028.4209, 1028.3718, 1028.3263, 1028.2704, 1028.214, 1028.1632, 1028.114, 1028.0631, 1028.0209, 1027.9728, 1027.9229, 1027.8784, 1027.8353, 1027.7915, 1027.7393, 1027.6866, 1027.6398, 1027.5863, 1027.536, 1027.4879, 1027.4331, 1027.3752, 1027.3157, 1027.2635, 1027.2112, 1027.1643, 1027.1093, 1027.0557, 1026.9841, 1026.9275, 1026.8313, 1026.7477, 1026.679, 1026.5774, 1026.4521, 1026.3759, 1026.2596, 1026.1709, 1026.0859, 1025.9141, 1025.7799, 1025.6495, 1025.4767, 1025.353, 1025.2007, 1025.0703, 1024.9423, 1024.8531, 1024.7645, 1024.6882, 1024.5398, 1024.2195, 1024.1619, NaN, NaN, 1029.277, 1029.2483, 1029.2133, 1029.1628, 1029.1146, 1029.0642, 1029.0149, 1028.963, 1028.9078, 1028.8513, 1028.8027, 1028.7537, 1028.7063, 1028.6514, 1028.5963, 1028.5404, 1028.4816, 1028.4286, 1028.3804, 1028.3374, 1028.2881, 1028.2344, 1028.1802, 1028.132, 1028.0787, 1028.0245, 1027.9756, 1027.922, 1027.8771, 1027.8282, 1027.7815, 1027.7261, 1027.6691, 1027.6149, 1027.5662, 1027.5067, 1027.4514, 1027.3993, 1027.3331, 1027.2778, 1027.2266, 1027.1759, 1027.1232, 1027.0497, 1026.9625, 1026.8627, 1026.7925, 1026.7218, 1026.6256, 1026.5334, 1026.4264, 1026.3073, 1026.2046, 1026.1102, 1026.0128, 1025.8977, 1025.6907, 1025.4729, 1025.3658, 1025.2579, 1025.0968, 1024.8947, 1024.7329, 1024.684, 1024.6378, 1024.6052, 1024.578, 1024.5686, NaN, NaN, 1029.2891, 1029.2612, 1029.2302, 1029.1835, 1029.1289, 1029.0763, 1029.0217, 1028.9749, 1028.9253, 1028.8726, 1028.8195, 1028.7709, 1028.718, 1028.6648, 1028.6125, 1028.5587, 1028.5071, 1028.4568, 1028.4064, 1028.3586, 1028.3086, 1028.2672, 1028.22, 1028.1698, 1028.1119, 1028.0519, 1028.0001, 1027.9535, 1027.9058, 1027.8513, 1027.8073, 1027.756, 1027.6992, 1027.6503, 1027.601, 1027.5482, 1027.4884, 1027.4329, 1027.3784, 1027.3264, 1027.2686, 1027.2136, 1027.1555, 1027.0797, 1027.0121, 1026.9388, 1026.8599, 1026.7959, 1026.6863, 1026.5989, 1026.5128, 1026.4011, 1026.2456, 1026.105, 1025.9824, 1025.8174, 1025.6346, 1025.5184, 1025.3909, 1025.2333, 1025.0482, 1024.7893, 1024.7087, 1024.6208, 1024.5323, 1024.4985, 1024.4684, 1024.4403, NaN, NaN, 1029.2792, 1029.252, 1029.2151, 1029.168, 1029.1147, 1029.0712, 1029.024, 1028.978, 1028.9325, 1028.885, 1028.8346, 1028.78, 1028.7345, 1028.685, 1028.6431, 1028.5929, 1028.5427, 1028.4977, 1028.4458, 1028.4039, 1028.3564, 1028.3071, 1028.2648, 1028.2158, 1028.1724, 1028.1294, 1028.0795, 1028.0306, 1027.9801, 1027.9255, 1027.875, 1027.8182, 1027.7659, 1027.7142, 1027.664, 1027.617, 1027.5691, 1027.515, 1027.4646, 1027.4125, 1027.3589, 1027.3002, 1027.2512, 1027.1974, 1027.1316, 1027.0822, 1027.027, 1026.9146, 1026.8223, 1026.7517, 1026.6584, 1026.5698, 1026.4778, 1026.3448, 1026.1844, 1026.0547, 1025.9153, 1025.75, 1025.6014, 1025.4321, 1025.2894, 1025.1962, 1025.0332, 1024.8312, 1024.6599, 1024.44, 1024.2759, 1024.1782, 1024.1473, 1024.1157, 1024.0891, NaN, NaN, 1029.2727, 1029.2385, 1029.2024, 1029.1588, 1029.107, 1029.0592, 1029.0154, 1028.9685, 1028.9264, 1028.8732, 1028.83, 1028.7878, 1028.7418, 1028.6923, 1028.6393, 1028.5906, 1028.5452, 1028.5039, 1028.4606, 1028.4149, 1028.369, 1028.3217, 1028.2712, 1028.2135, 1028.164, 1028.1144, 1028.0653, 1028.0227, 1027.9741, 1027.9193, 1027.873, 1027.8273, 1027.7788, 1027.7311, 1027.6906, 1027.6433, 1027.5951, 1027.5492, 1027.5005, 1027.4515, 1027.4027, 1027.3513, 1027.2925, 1027.2367, 1027.1848, 1027.1426, 1027.0731, 1026.991, 1026.911, 1026.8007, 1026.7126, 1026.6648, 1026.5737, 1026.4722, 1026.3174, 1026.0941, 1025.9359, 1025.8279, 1025.7253, 1025.6298, 1025.5033, 1025.396, 1025.2782, 1025.1857, 1025.0304, 1024.8696, 1024.7738, 1024.7046, 1024.5978, 1024.4724, 1024.2101, 1024.0452, NaN, NaN, 1029.2736, 1029.2427, 1029.1993, 1029.1539, 1029.1036, 1029.055, 1029.0057, 1028.9647, 1028.92, 1028.8718, 1028.8201, 1028.7633, 1028.7125, 1028.6643, 1028.615, 1028.5674, 1028.5162, 1028.4657, 1028.4174, 1028.3699, 1028.3203, 1028.2657, 1028.2126, 1028.1624, 1028.1042, 1028.0549, 1028.0016, 1027.9496, 1027.9008, 1027.8513, 1027.8015, 1027.7484, 1027.7026, 1027.66, 1027.6053, 1027.5513, 1027.4984, 1027.4485, 1027.3942, 1027.3401, 1027.2904, 1027.2316, 1027.1641, 1027.1084, 1027.0735, 1027.0186, 1026.9221, 1026.8138, 1026.732, 1026.658, 1026.5964, 1026.5366, 1026.4445, 1026.3682, 1026.2686, 1026.177, 1026.0995, 1026.027, 1025.918, 1025.8401, 1025.7535, 1025.6198, 1025.4679, 1025.3529, 1025.2589, 1025.1184, 1025.0358, 1024.9324, 1024.8278, 1024.7555, 1024.6984, 1024.6332, 1024.4775, 1024.2057, 1024.165, NaN, NaN, 1029.2921, 1029.2635, 1029.2284, 1029.1869, 1029.1368, 1029.0841, 1029.0319, 1028.9811, 1028.9341, 1028.8854, 1028.8442, 1028.799, 1028.7416, 1028.6866, 1028.6372, 1028.5896, 1028.5464, 1028.4985, 1028.4437, 1028.4042, 1028.361, 1028.31, 1028.2601, 1028.2162, 1028.164, 1028.1167, 1028.071, 1028.0208, 1027.9747, 1027.9221, 1027.8708, 1027.8164, 1027.764, 1027.7148, 1027.649, 1027.5986, 1027.5469, 1027.4951, 1027.4517, 1027.3934, 1027.3298, 1027.274, 1027.2133, 1027.1606, 1027.1144, 1027.0573, 1026.9941, 1026.9319, 1026.868, 1026.7607, 1026.626, 1026.5597, 1026.4547, 1026.355, 1026.2178, 1026.097, 1025.9556, 1025.8352, 1025.6854, 1025.5566, 1025.4099, 1025.2168, 1025.0778, 1024.9269, 1024.7432, 1024.6976, 1024.637, 1024.4551, 1024.3112, NaN, NaN, 1029.2911, 1029.264, 1029.2268, 1029.1744, 1029.1215, 1029.0775, 1029.0281, 1028.9746, 1028.9264, 1028.874, 1028.8297, 1028.7798, 1028.709, 1028.6553, 1028.6058, 1028.5524, 1028.5013, 1028.4501, 1028.3973, 1028.3442, 1028.2952, 1028.2439, 1028.1942, 1028.141, 1028.0869, 1028.0334, 1027.9797, 1027.9268, 1027.8796, 1027.8331, 1027.7872, 1027.7289, 1027.6699, 1027.6171, 1027.5724, 1027.5269, 1027.4685, 1027.4192, 1027.3698, 1027.3174, 1027.2695, 1027.2156, 1027.1644, 1027.1168, 1027.0549, 1026.9916, 1026.9152, 1026.813, 1026.6864, 1026.6135, 1026.5342, 1026.4392, 1026.2947, 1026.1364, 1025.9584, 1025.8141, 1025.6431, 1025.47, 1025.3424, 1025.2307, 1025.1184, 1024.9955, 1024.8889, 1024.8022, 1024.6956, 1024.5818, 1024.4589, 1024.4437, NaN, NaN, 1029.2788, 1029.2512, 1029.2158, 1029.1598, 1029.1091, 1029.0505, 1028.995, 1028.9509, 1028.9006, 1028.8457, 1028.7982, 1028.7418, 1028.6932, 1028.6417, 1028.5952, 1028.5487, 1028.5002, 1028.4525, 1028.4072, 1028.3566, 1028.3082, 1028.2563, 1028.199, 1028.1499, 1028.0907, 1028.034, 1027.9884, 1027.9391, 1027.8915, 1027.8398, 1027.7858, 1027.7317, 1027.6836, 1027.6329, 1027.5757, 1027.5232, 1027.4749, 1027.4258, 1027.3768, 1027.3258, 1027.2661, 1027.2075, 1027.1608, 1027.108, 1027.054, 1026.9681, 1026.9008, 1026.8151, 1026.723, 1026.6495, 1026.566, 1026.4298, 1026.267, 1026.1155, 1025.9747, 1025.8755, 1025.7975, 1025.6809, 1025.5051, 1025.3755, 1025.2245, 1025.1023, 1025.0092, 1024.8159, 1024.7358, 1024.6946, 1024.6498, 1024.5642, 1024.3423, 1024.2325, NaN, NaN, 1029.2688, 1029.2424, 1029.2015, 1029.1482, 1029.0927, 1029.0374, 1028.9894, 1028.9473, 1028.8953, 1028.8461, 1028.7991, 1028.7465, 1028.6942, 1028.6478, 1028.5948, 1028.5448, 1028.497, 1028.445, 1028.3915, 1028.337, 1028.2803, 1028.2281, 1028.1783, 1028.1276, 1028.0751, 1028.0186, 1027.9717, 1027.9233, 1027.87, 1027.819, 1027.7759, 1027.7234, 1027.667, 1027.6177, 1027.5712, 1027.5265, 1027.4773, 1027.416, 1027.3561, 1027.2997, 1027.2512, 1027.1982, 1027.1464, 1027.0854, 1027.0266, 1026.9537, 1026.8854, 1026.7908, 1026.6802, 1026.6191, 1026.5144, 1026.4133, 1026.288, 1026.1758, 1026.0479, 1025.9628, 1025.848, 1025.7054, 1025.4766, 1025.3553, 1025.1746, 1024.9974, 1024.8685, 1024.697, 1024.4377, 1024.1414, 1024.103, 1024.0906, NaN, NaN, 1029.2701, 1029.2388, 1029.201, 1029.1483, 1029.1025, 1029.0487, 1029.0042, 1028.9546, 1028.9047, 1028.8552, 1028.803, 1028.7489, 1028.7043, 1028.6613, 1028.6138, 1028.5637, 1028.5126, 1028.4578, 1028.4133, 1028.3661, 1028.3188, 1028.2726, 1028.2233, 1028.1768, 1028.1237, 1028.074, 1028.0243, 1027.9802, 1027.929, 1027.8739, 1027.8215, 1027.7635, 1027.7064, 1027.6653, 1027.6234, 1027.5681, 1027.5082, 1027.4589, 1027.3993, 1027.3376, 1027.287, 1027.2402, 1027.171, 1027.1115, 1027.0529, 1026.9982, 1026.9193, 1026.8545, 1026.7339, 1026.6288, 1026.5284, 1026.441, 1026.3431, 1026.2235, 1026.0675, 1025.9624, 1025.8658, 1025.7448, 1025.5929, 1025.4364, 1025.3282, 1025.1738, 1024.9895, 1024.8795, 1024.7488, 1024.581, 1024.3281, 1024.2068, NaN, NaN, 1029.2976, 1029.2686, 1029.2286, 1029.1769, 1029.1257, 1029.0724, 1029.0251, 1028.9749, 1028.9282, 1028.8774, 1028.8268, 1028.7806, 1028.7307, 1028.6829, 1028.6394, 1028.5933, 1028.5435, 1028.4894, 1028.4419, 1028.3938, 1028.3427, 1028.2942, 1028.247, 1028.1973, 1028.1509, 1028.1013, 1028.053, 1028.0094, 1027.9608, 1027.9103, 1027.8646, 1027.8119, 1027.7607, 1027.7129, 1027.6632, 1027.6195, 1027.5657, 1027.5015, 1027.4427, 1027.3934, 1027.338, 1027.2765, 1027.2137, 1027.1643, 1027.1089, 1027.0543, 1026.9844, 1026.9229, 1026.835, 1026.7504, 1026.6924, 1026.6067, 1026.4977, 1026.4103, 1026.3142, 1026.2029, 1026.0612, 1025.9652, 1025.8021, 1025.6886, 1025.4972, 1025.2854, 1025.1359, 1024.9143, 1024.8086, 1024.761, 1024.7163, 1024.6289, 1024.4784, 1024.3164, 1024.2979, NaN, NaN, 1029.29, 1029.2634, 1029.2302, 1029.1815, 1029.1339, 1029.0776, 1029.0238, 1028.972, 1028.9197, 1028.8693, 1028.8273, 1028.7769, 1028.7272, 1028.6837, 1028.6368, 1028.589, 1028.5366, 1028.4874, 1028.4381, 1028.394, 1028.3416, 1028.2894, 1028.2423, 1028.1924, 1028.1459, 1028.0972, 1028.0461, 1027.9926, 1027.9452, 1027.8917, 1027.8427, 1027.7828, 1027.7239, 1027.672, 1027.6145, 1027.5615, 1027.4923, 1027.4193, 1027.3495, 1027.2963, 1027.2314, 1027.1699, 1027.0984, 1027.0339, 1026.9742, 1026.8777, 1026.7585, 1026.6915, 1026.574, 1026.4266, 1026.2623, 1026.0671, 1025.9486, 1025.7856, 1025.6879, 1025.5134, 1025.3857, 1025.3098, 1025.1908, 1025.0916, 1024.9639, 1024.7651, 1024.7052, 1024.5059, 1024.4225, 1024.2653, 1024.1633, NaN, NaN, 1029.2858, 1029.2567, 1029.2203, 1029.1696, 1029.1187, 1029.0665, 1029.0183, 1028.9711, 1028.9258, 1028.8801, 1028.835, 1028.7908, 1028.7396, 1028.6918, 1028.6449, 1028.5974, 1028.5394, 1028.4912, 1028.4424, 1028.3893, 1028.3408, 1028.2822, 1028.2307, 1028.1765, 1028.1284, 1028.077, 1028.0243, 1027.9716, 1027.9127, 1027.8618, 1027.8015, 1027.7555, 1027.7068, 1027.6492, 1027.5996, 1027.5555, 1027.4991, 1027.4397, 1027.3832, 1027.336, 1027.2822, 1027.2201, 1027.1599, 1027.0988, 1027.0295, 1026.9446, 1026.8553, 1026.7845, 1026.7092, 1026.5881, 1026.4932, 1026.3425, 1026.1694, 1026.0658, 1025.9559, 1025.8077, 1025.7079, 1025.652, 1025.5498, 1025.4109, 1025.295, 1025.1182, 1024.9742, 1024.873, 1024.7516, 1024.6387, 1024.5316, 1024.4207, NaN, NaN, 1029.2604, 1029.2351, 1029.1956, 1029.146, 1029.0994, 1029.0471, 1028.9933, 1028.9397, 1028.8938, 1028.8442, 1028.7968, 1028.7478, 1028.698, 1028.6411, 1028.5911, 1028.539, 1028.4875, 1028.4259, 1028.3701, 1028.3164, 1028.2662, 1028.2158, 1028.1658, 1028.1124, 1028.0599, 1028.0094, 1027.9573, 1027.9026, 1027.8451, 1027.8011, 1027.7515, 1027.7034, 1027.6598, 1027.6068, 1027.5508, 1027.5015, 1027.451, 1027.4037, 1027.3446, 1027.2786, 1027.2053, 1027.1584, 1027.1096, 1027.0416, 1026.9855, 1026.9178, 1026.8387, 1026.747, 1026.6486, 1026.5519, 1026.4453, 1026.3475, 1026.2328, 1026.1256, 1026.0541, 1025.8716, 1025.7177, 1025.5907, 1025.4734, 1025.358, 1025.2819, 1025.1195, 1025.046, 1024.9558, 1024.8209, 1024.6023, 1024.5051, 1024.2983, 1024.2312, NaN, NaN, 1029.2799, 1029.2544, 1029.2206, 1029.1748, 1029.1259, 1029.0754, 1029.0245, 1028.9692, 1028.9214, 1028.873, 1028.8228, 1028.7697, 1028.7155, 1028.6626, 1028.6125, 1028.5642, 1028.5177, 1028.4707, 1028.4219, 1028.3622, 1028.3119, 1028.2626, 1028.2114, 1028.1555, 1028.1033, 1028.0529, 1027.9998, 1027.9478, 1027.8862, 1027.8314, 1027.7869, 1027.7383, 1027.6814, 1027.6282, 1027.5815, 1027.5282, 1027.4747, 1027.42, 1027.3582, 1027.3035, 1027.2356, 1027.167, 1027.1122, 1027.0519, 1026.9845, 1026.9069, 1026.8204, 1026.7264, 1026.6533, 1026.55, 1026.4794, 1026.385, 1026.2677, 1026.171, 1026.0394, 1025.833, 1025.7161, 1025.5757, 1025.4255, 1025.2607, 1025.159, 1025.0054, 1024.8866, 1024.772, 1024.6829, 1024.646, 1024.6093, 1024.5619, 1024.5457, NaN, NaN, 1029.2659, 1029.239, 1029.2004, 1029.1506, 1029.097, 1029.0508, 1029.0035, 1028.9518, 1028.9065, 1028.8643, 1028.8186, 1028.7728, 1028.7272, 1028.6824, 1028.6339, 1028.5912, 1028.5455, 1028.4998, 1028.4514, 1028.3961, 1028.3441, 1028.2985, 1028.2549, 1028.205, 1028.1578, 1028.1105, 1028.065, 1028.0183, 1027.9757, 1027.929, 1027.8809, 1027.8345, 1027.7892, 1027.731, 1027.6792, 1027.6304, 1027.5925, 1027.5428, 1027.4946, 1027.439, 1027.3918, 1027.3242, 1027.2754, 1027.2197, 1027.1525, 1027.102, 1027.0426, 1026.9766, 1026.9054, 1026.8374, 1026.761, 1026.6611, 1026.5358, 1026.4353, 1026.3152, 1026.1995, 1026.0438, 1025.8743, 1025.7114, 1025.5355, 1025.45, 1025.346, 1025.0726, 1024.9309, 1024.8754, 1024.7872, 1024.6976, 1024.6698, 1024.6501, 1024.6276, 1024.6023, 1024.58, NaN, NaN, 1029.2877, 1029.2579, 1029.2205, 1029.1697, 1029.1213, 1029.0737, 1029.02, 1028.9722, 1028.9292, 1028.8834, 1028.8362, 1028.7861, 1028.7294, 1028.681, 1028.6335, 1028.5856, 1028.5331, 1028.4855, 1028.4305, 1028.3744, 1028.3204, 1028.2697, 1028.2263, 1028.1781, 1028.1278, 1028.0748, 1028.022, 1027.974, 1027.9297, 1027.8763, 1027.8235, 1027.7771, 1027.7316, 1027.6864, 1027.6355, 1027.5817, 1027.5405, 1027.4917, 1027.4429, 1027.3864, 1027.3279, 1027.2731, 1027.2106, 1027.1543, 1027.0803, 1027.013, 1026.9457, 1026.86, 1026.7523, 1026.6404, 1026.5424, 1026.4313, 1026.287, 1026.1577, 1026.0262, 1025.8885, 1025.7749, 1025.6251, 1025.5505, 1025.4258, 1025.2793, 1025.1671, 1024.8915, 1024.7134, 1024.5906, 1024.497, 1024.3423, 1024.2277, 1024.2094, NaN, NaN, 1029.2771, 1029.2483, 1029.2128, 1029.1646, 1029.1188, 1029.0688, 1029.0194, 1028.9739, 1028.9292, 1028.8839, 1028.8356, 1028.7903, 1028.7463, 1028.703, 1028.6617, 1028.6252, 1028.5815, 1028.5344, 1028.4922, 1028.438, 1028.3843, 1028.3359, 1028.2821, 1028.23, 1028.1727, 1028.1183, 1028.0577, 1027.9983, 1027.9419, 1027.8895, 1027.841, 1027.7872, 1027.7365, 1027.6874, 1027.6335, 1027.5875, 1027.5364, 1027.4874, 1027.4436, 1027.392, 1027.3253, 1027.2775, 1027.2085, 1027.1401, 1027.0829, 1027.0033, 1026.9421, 1026.8667, 1026.7716, 1026.6804, 1026.5906, 1026.5115, 1026.4076, 1026.2545, 1026.1462, 1026.0052, 1025.8767, 1025.7577, 1025.6605, 1025.5883, 1025.5057, 1025.402, 1025.3147, 1025.1593, 1024.9645, 1024.8336, 1024.6254, 1024.4291, 1024.3607, 1024.2365, 1024.1946, 1024.1832, NaN, NaN, 1029.2853, 1029.26, 1029.2247, 1029.1708, 1029.1161, 1029.0668, 1029.0144, 1028.9584, 1028.9044, 1028.853, 1028.8029, 1028.7493, 1028.6981, 1028.6492, 1028.5991, 1028.5474, 1028.4952, 1028.4436, 1028.3894, 1028.335, 1028.2788, 1028.2327, 1028.1819, 1028.1367, 1028.0817, 1028.0223, 1027.9789, 1027.9309, 1027.8846, 1027.8364, 1027.7842, 1027.7241, 1027.6746, 1027.6246, 1027.5693, 1027.5228, 1027.4755, 1027.4292, 1027.3839, 1027.3406, 1027.2837, 1027.2279, 1027.1569, 1027.0972, 1027.0564, 1026.9778, 1026.9137, 1026.8499, 1026.7827, 1026.7162, 1026.6007, 1026.5009, 1026.378, 1026.197, 1026.0845, 1025.9487, 1025.8042, 1025.6136, 1025.5056, 1025.3743, 1025.2499, 1025.0968, 1024.9763, 1024.8121, 1024.6389, 1024.5873, 1024.542, 1024.4545, 1024.3898, NaN, NaN, 1029.2837, 1029.2528, 1029.2158, 1029.1675, 1029.1136, 1029.0607, 1029.0103, 1028.9614, 1028.9138, 1028.8611, 1028.8171, 1028.7709, 1028.722, 1028.6687, 1028.6193, 1028.5747, 1028.5262, 1028.4802, 1028.4309, 1028.3829, 1028.3309, 1028.2773, 1028.225, 1028.1708, 1028.1208, 1028.0654, 1028.0195, 1027.9683, 1027.9121, 1027.8667, 1027.8203, 1027.7643, 1027.7041, 1027.6482, 1027.5963, 1027.5367, 1027.472, 1027.4177, 1027.3652, 1027.3079, 1027.2529, 1027.208, 1027.1431, 1027.0645, 1027.0107, 1026.9495, 1026.8691, 1026.7883, 1026.6969, 1026.599, 1026.4971, 1026.4059, 1026.2428, 1026.1069, 1025.9883, 1025.7938, 1025.6234, 1025.4828, 1025.3667, 1025.27, 1025.1033, 1024.9917, 1024.8738, 1024.6573, 1024.4894, 1024.4146, 1024.3147, 1024.2719, NaN, NaN, 1029.284, 1029.2568, 1029.2225, 1029.1713, 1029.1222, 1029.0695, 1029.0195, 1028.9668, 1028.9147, 1028.8661, 1028.8126, 1028.7654, 1028.7137, 1028.6686, 1028.6246, 1028.5771, 1028.5344, 1028.4889, 1028.4434, 1028.3942, 1028.3434, 1028.2997, 1028.2563, 1028.2114, 1028.158, 1028.1082, 1028.0671, 1028.0193, 1027.971, 1027.9258, 1027.8733, 1027.8247, 1027.7756, 1027.7183, 1027.6711, 1027.6166, 1027.5485, 1027.4956, 1027.429, 1027.3737, 1027.3184, 1027.2538, 1027.2052, 1027.1454, 1027.0789, 1026.9952, 1026.8872, 1026.8011, 1026.7086, 1026.597, 1026.4609, 1026.2979, 1026.1724, 1026.0088, 1025.8785, 1025.7335, 1025.5885, 1025.4982, 1025.3549, 1025.2428, 1025.182, 1025.0851, 1024.9468, 1024.8086, 1024.7617, 1024.696, 1024.6444, 1024.5844, 1024.5562, NaN, NaN, 1029.2955, 1029.2694, 1029.2356, 1029.1885, 1029.1436, 1029.1003, 1029.0514, 1029.0026, 1028.954, 1028.9086, 1028.8661, 1028.8185, 1028.7694, 1028.7185, 1028.6665, 1028.6151, 1028.5603, 1028.5061, 1028.4521, 1028.4033, 1028.3433, 1028.2935, 1028.2448, 1028.1915, 1028.1436, 1028.084, 1028.0328, 1027.9763, 1027.9277, 1027.8856, 1027.8342, 1027.7809, 1027.7316, 1027.6844, 1027.632, 1027.5796, 1027.5209, 1027.4631, 1027.407, 1027.3634, 1027.3043, 1027.242, 1027.173, 1027.1058, 1027.0327, 1026.9586, 1026.8914, 1026.8091, 1026.7318, 1026.6316, 1026.5123, 1026.3435, 1026.2297, 1026.0962, 1025.952, 1025.8456, 1025.7378, 1025.5963, 1025.5132, 1025.3896, 1025.3016, 1025.1875, 1025.0315, 1024.8749, 1024.7753, 1024.6722, 1024.6263, 1024.5956, 1024.5812, NaN, NaN, 1029.2568, 1029.2274, 1029.1918, 1029.1492, 1029.1079, 1029.0619, 1029.0159, 1028.969, 1028.9233, 1028.8779, 1028.8269, 1028.7828, 1028.7365, 1028.6925, 1028.6454, 1028.5967, 1028.5453, 1028.4968, 1028.4482, 1028.3961, 1028.3468, 1028.2947, 1028.2395, 1028.1836, 1028.1329, 1028.0808, 1028.0271, 1027.9764, 1027.922, 1027.8676, 1027.8181, 1027.7728, 1027.7228, 1027.6702, 1027.6229, 1027.5691, 1027.5089, 1027.4546, 1027.4055, 1027.3516, 1027.2916, 1027.2231, 1027.1337, 1027.0741, 1027.0244, 1026.9666, 1026.9022, 1026.8206, 1026.7308, 1026.6172, 1026.5037, 1026.3816, 1026.2344, 1026.0912, 1025.9646, 1025.8458, 1025.6711, 1025.5457, 1025.4414, 1025.3099, 1025.1188, 1024.9021, 1024.8271, 1024.7068, 1024.6417, 1024.6108, 1024.5818, 1024.562, NaN, NaN, 1029.2892, 1029.259, 1029.2236, 1029.1754, 1029.1328, 1029.0837, 1029.0369, 1028.9866, 1028.9379, 1028.8894, 1028.8428, 1028.7921, 1028.7401, 1028.6932, 1028.6447, 1028.5975, 1028.549, 1028.5001, 1028.4474, 1028.3984, 1028.3483, 1028.2933, 1028.2415, 1028.1915, 1028.1394, 1028.0757, 1028.0254, 1027.9741, 1027.9221, 1027.8706, 1027.8207, 1027.7694, 1027.7144, 1027.6674, 1027.6171, 1027.5625, 1027.509, 1027.4517, 1027.4015, 1027.3425, 1027.2902, 1027.2268, 1027.1575, 1027.1144, 1027.0509, 1026.995, 1026.9038, 1026.8556, 1026.7408, 1026.6558, 1026.5452, 1026.4222, 1026.2607, 1026.1329, 1026.0046, 1025.8438, 1025.7185, 1025.5894, 1025.4766, 1025.2238, 1025.0485, 1024.9113, 1024.847, 1024.7767, 1024.657, 1024.5845, 1024.5422, 1024.5139, 1024.4958, NaN, NaN, 1029.2776, 1029.2474, 1029.2057, 1029.1595, 1029.1075, 1029.0505, 1028.9943, 1028.9381, 1028.8821, 1028.8356, 1028.7828, 1028.7317, 1028.6826, 1028.6307, 1028.5789, 1028.5267, 1028.4762, 1028.4252, 1028.37, 1028.3151, 1028.2556, 1028.2032, 1028.1454, 1028.0895, 1028.0344, 1027.9792, 1027.9187, 1027.8647, 1027.8083, 1027.749, 1027.6907, 1027.6289, 1027.5701, 1027.5122, 1027.4634, 1027.4069, 1027.3524, 1027.293, 1027.2314, 1027.1793, 1027.1064, 1027.0284, 1026.9633, 1026.8873, 1026.8231, 1026.7488, 1026.6516, 1026.5564, 1026.4557, 1026.2694, 1026.1357, 1026.0168, 1025.8801, 1025.7345, 1025.616, 1025.4691, 1025.2776, 1025.1658, 1025.0199, 1024.8517, 1024.781, 1024.697, 1024.629, 1024.567, 1024.5227, 1024.4994, NaN, NaN, 1029.2815, 1029.2546, 1029.2214, 1029.1719, 1029.1185, 1029.0643, 1029.0133, 1028.9634, 1028.9158, 1028.8699, 1028.8204, 1028.7719, 1028.721, 1028.6737, 1028.6283, 1028.5837, 1028.5348, 1028.4927, 1028.447, 1028.3978, 1028.35, 1028.3085, 1028.26, 1028.2144, 1028.1671, 1028.1201, 1028.0706, 1028.0204, 1027.9763, 1027.9296, 1027.8716, 1027.8206, 1027.7705, 1027.7147, 1027.6604, 1027.5994, 1027.5455, 1027.489, 1027.437, 1027.3844, 1027.3153, 1027.2505, 1027.1718, 1027.0939, 1027.0416, 1026.9819, 1026.9115, 1026.8245, 1026.7351, 1026.6613, 1026.5698, 1026.454, 1026.3048, 1026.1781, 1026.069, 1025.9678, 1025.8336, 1025.68, 1025.5302, 1025.4049, 1025.243, 1025.074, 1024.8999, 1024.7421, 1024.5892, 1024.538, 1024.4733, 1024.4336, 1024.4055, 1024.374, 1024.3593, NaN, NaN, 1029.2573, 1029.2296, 1029.1917, 1029.1448, 1029.0906, 1029.0371, 1028.9857, 1028.9308, 1028.8827, 1028.8319, 1028.784, 1028.737, 1028.6919, 1028.6482, 1028.6001, 1028.5542, 1028.5012, 1028.4531, 1028.4025, 1028.3558, 1028.3053, 1028.2467, 1028.1976, 1028.1514, 1028.1006, 1028.054, 1028.0076, 1027.962, 1027.9064, 1027.8506, 1027.7933, 1027.7402, 1027.6918, 1027.6348, 1027.581, 1027.5256, 1027.4702, 1027.4111, 1027.3458, 1027.2832, 1027.2112, 1027.153, 1027.0995, 1027.0359, 1026.9584, 1026.8765, 1026.775, 1026.6981, 1026.592, 1026.476, 1026.3556, 1026.2612, 1026.1315, 1026.004, 1025.8431, 1025.6927, 1025.5594, 1025.4738, 1025.352, 1025.2356, 1025.1196, 1025.0093, 1024.8157, 1024.5724, 1024.3722, 1024.3411, 1024.3099, 1024.2578, 1024.1978, 1024.1705, NaN, NaN, 1029.2693, 1029.2395, 1029.2025, 1029.1493, 1029.0979, 1029.0457, 1028.9935, 1028.9392, 1028.8835, 1028.8344, 1028.7819, 1028.7356, 1028.6906, 1028.6365, 1028.5814, 1028.5374, 1028.4889, 1028.4425, 1028.3911, 1028.3387, 1028.293, 1028.2463, 1028.2002, 1028.1593, 1028.1075, 1028.054, 1027.9983, 1027.9463, 1027.8923, 1027.8384, 1027.7823, 1027.7303, 1027.6825, 1027.6288, 1027.5774, 1027.5221, 1027.4739, 1027.4204, 1027.3635, 1027.3091, 1027.2501, 1027.1705, 1027.1146, 1027.0465, 1026.9961, 1026.9264, 1026.8574, 1026.7726, 1026.6842, 1026.5663, 1026.4529, 1026.3398, 1026.1835, 1026.0215, 1025.9077, 1025.7831, 1025.6437, 1025.5354, 1025.3954, 1025.255, 1025.0923, 1024.9624, 1024.7153, 1024.4587, 1024.328, 1024.2639, 1024.2045, 1024.1635, 1024.1456, NaN, NaN, 1029.2594, 1029.2302, 1029.1942, 1029.1427, 1029.0812, 1029.0277, 1028.9739, 1028.9203, 1028.8696, 1028.8136, 1028.7625, 1028.708, 1028.6556, 1028.6027, 1028.5479, 1028.489, 1028.4386, 1028.3898, 1028.3412, 1028.295, 1028.244, 1028.1921, 1028.1378, 1028.0853, 1028.0306, 1027.9741, 1027.9229, 1027.8713, 1027.8179, 1027.756, 1027.7141, 1027.6731, 1027.6187, 1027.5675, 1027.5204, 1027.4617, 1027.4, 1027.3407, 1027.2821, 1027.2168, 1027.166, 1027.0906, 1027.0135, 1026.9253, 1026.8403, 1026.7578, 1026.6752, 1026.5626, 1026.47, 1026.3607, 1026.2141, 1026.0582, 1025.9083, 1025.727, 1025.5968, 1025.4458, 1025.313, 1025.1971, 1025.0868, 1024.9706, 1024.8474, 1024.6731, 1024.4281, 1024.364, 1024.34, 1024.3079, 1024.252, 1024.2135, 1024.1946, NaN, NaN, 1029.2892, 1029.2611, 1029.2246, 1029.1703, 1029.1256, 1029.0798, 1029.0344, 1028.9875, 1028.9421, 1028.8988, 1028.8516, 1028.8015, 1028.7562, 1028.7086, 1028.6592, 1028.6113, 1028.564, 1028.5184, 1028.468, 1028.4186, 1028.3733, 1028.3279, 1028.2808, 1028.2343, 1028.1805, 1028.1382, 1028.0887, 1028.0345, 1027.9856, 1027.9329, 1027.8816, 1027.8334, 1027.7872, 1027.7422, 1027.6995, 1027.6527, 1027.6041, 1027.555, 1027.5073, 1027.459, 1027.4072, 1027.3552, 1027.2979, 1027.237, 1027.1731, 1027.1053, 1027.0216, 1026.9347, 1026.8575, 1026.7565, 1026.6312, 1026.5121, 1026.3945, 1026.2622, 1026.1316, 1025.9961, 1025.8126, 1025.7294, 1025.6102, 1025.4543, 1025.3416, 1025.2568, 1025.1365, 1025.0605, 1024.9592, 1024.8425, 1024.6582, 1024.4562, 1024.2808, 1024.251, 1024.2179, 1024.1951, 1024.1573, 1024.117, NaN, NaN, 1029.2734, 1029.246, 1029.2094, 1029.1595, 1029.1058, 1029.0491, 1028.9965, 1028.9452, 1028.8934, 1028.8412, 1028.7886, 1028.7363, 1028.6829, 1028.6342, 1028.587, 1028.5427, 1028.4926, 1028.4412, 1028.395, 1028.35, 1028.3016, 1028.2529, 1028.2031, 1028.1522, 1028.1062, 1028.0586, 1028.0082, 1027.9553, 1027.9045, 1027.8583, 1027.8108, 1027.7637, 1027.7008, 1027.6459, 1027.5912, 1027.5382, 1027.4899, 1027.4368, 1027.3784, 1027.3091, 1027.248, 1027.1993, 1027.1407, 1027.0485, 1026.9518, 1026.8724, 1026.8027, 1026.7003, 1026.6302, 1026.537, 1026.4441, 1026.2844, 1026.1511, 1026.0001, 1025.8254, 1025.673, 1025.5515, 1025.4459, 1025.3007, 1025.1571, 1025.0692, 1025.0052, 1024.8468, 1024.681, 1024.4023, 1024.2288, 1024.2019, 1024.1758, 1024.1482, 1024.1188, 1024.0787, NaN, NaN, 1029.2554, 1029.2295, 1029.1951, 1029.1466, 1029.0964, 1029.0482, 1029.0022, 1028.9537, 1028.9049, 1028.8549, 1028.8025, 1028.7554, 1028.709, 1028.6609, 1028.6116, 1028.5671, 1028.5104, 1028.457, 1028.4032, 1028.3507, 1028.297, 1028.2511, 1028.2003, 1028.1458, 1028.0901, 1028.0374, 1027.9921, 1027.9392, 1027.8887, 1027.8372, 1027.7833, 1027.7333, 1027.6841, 1027.629, 1027.5773, 1027.5253, 1027.4697, 1027.4156, 1027.3517, 1027.2887, 1027.2229, 1027.1624, 1027.0962, 1027.0402, 1026.9622, 1026.8679, 1026.7621, 1026.6708, 1026.5894, 1026.4971, 1026.3646, 1026.1995, 1026.0397, 1025.9178, 1025.8212, 1025.6932, 1025.5498, 1025.4081, 1025.2351, 1025.1616, 1025.0717, 1024.9546, 1024.8652, 1024.6614, 1024.3087, 1024.2389, 1024.1998, 1024.1561, 1024.1079, 1024.0288, 1023.9432, 1023.9223, NaN, NaN, 1029.2333, 1029.2074, 1029.1768, 1029.1346, 1029.092, 1029.0533, 1029.0098, 1028.9645, 1028.9242, 1028.8832, 1028.8383, 1028.793, 1028.7477, 1028.7017, 1028.6516, 1028.6064, 1028.5598, 1028.5165, 1028.4694, 1028.4213, 1028.3761, 1028.3301, 1028.2845, 1028.2415, 1028.1941, 1028.151, 1028.105, 1028.0583, 1028.0094, 1027.9628, 1027.9147, 1027.868, 1027.8215, 1027.7732, 1027.7252, 1027.6813, 1027.6321, 1027.5879, 1027.5394, 1027.49, 1027.4432, 1027.3998, 1027.3491, 1027.3019, 1027.2396, 1027.1674, 1027.0968, 1027.0404, 1026.965, 1026.8832, 1026.8069, 1026.7274, 1026.6313, 1026.508, 1026.3805, 1026.2728, 1026.1351, 1026.0157, 1025.8513, 1025.7568, 1025.5717, 1025.4359, 1025.3279, 1025.1937, 1025.1263, 1025.0084, 1024.8551, 1024.769, 1024.5702, 1024.3096, 1024.1189, 1024.0225, 1024.0011, 1023.97943, 1023.9521, 1023.92413, 1023.9043, NaN, NaN, 1029.2626, 1029.233, 1029.198, 1029.1514, 1029.0995, 1029.0452, 1028.9965, 1028.9443, 1028.893, 1028.8386, 1028.7896, 1028.7343, 1028.6735, 1028.6147, 1028.5588, 1028.5043, 1028.4537, 1028.4032, 1028.347, 1028.293, 1028.2428, 1028.1946, 1028.1444, 1028.0925, 1028.0441, 1027.9907, 1027.9376, 1027.8807, 1027.8285, 1027.7827, 1027.7362, 1027.6832, 1027.6133, 1027.5524, 1027.4934, 1027.4266, 1027.3556, 1027.2887, 1027.2296, 1027.1641, 1027.0972, 1027.0131, 1026.9379, 1026.85, 1026.7582, 1026.6355, 1026.5103, 1026.423, 1026.265, 1026.0817, 1025.9001, 1025.7633, 1025.6431, 1025.5476, 1025.4303, 1025.3193, 1025.2335, 1025.1201, 1025.0251, 1024.9121, 1024.8114, 1024.675, 1024.4169, 1024.1599, 1024.0425, 1024.0034, 1023.977, 1023.9529, 1023.93134, 1023.9175, NaN, NaN, 1029.2571, 1029.2311, 1029.1993, 1029.148, 1029.0963, 1029.0426, 1028.9946, 1028.9427, 1028.8969, 1028.8453, 1028.7965, 1028.7457, 1028.6979, 1028.6454, 1028.5918, 1028.5416, 1028.4923, 1028.4362, 1028.3856, 1028.3389, 1028.2906, 1028.2439, 1028.1997, 1028.1538, 1028.1099, 1028.0602, 1028.0134, 1027.9596, 1027.91, 1027.8575, 1027.8009, 1027.754, 1027.7087, 1027.6588, 1027.6062, 1027.5474, 1027.4968, 1027.4402, 1027.3826, 1027.3174, 1027.2695, 1027.1993, 1027.1135, 1027.0552, 1026.986, 1026.8997, 1026.8247, 1026.724, 1026.6215, 1026.4976, 1026.3416, 1026.2239, 1026.1045, 1025.9562, 1025.8164, 1025.6788, 1025.5659, 1025.4979, 1025.3708, 1025.2618, 1025.1417, 1025.08, 1024.9924, 1024.8622, 1024.5697, 1024.3387, 1024.165, 1024.066, 1024.0378, 1024.0166, 1023.9943, 1023.9709, 1023.9463, NaN, NaN, 1029.2637, 1029.2413, 1029.2067, 1029.162, 1029.116, 1029.0673, 1029.0146, 1028.966, 1028.9155, 1028.8661, 1028.8171, 1028.7664, 1028.7112, 1028.6604, 1028.6057, 1028.5546, 1028.5043, 1028.4471, 1028.3894, 1028.3271, 1028.2684, 1028.2146, 1028.1704, 1028.1202, 1028.0767, 1028.0333, 1027.9819, 1027.9248, 1027.8717, 1027.816, 1027.7627, 1027.7119, 1027.6675, 1027.6062, 1027.5591, 1027.4926, 1027.4255, 1027.3694, 1027.3251, 1027.2725, 1027.2085, 1027.1381, 1027.0631, 1026.99, 1026.9121, 1026.8251, 1026.7406, 1026.6147, 1026.5111, 1026.3405, 1026.1603, 1025.9962, 1025.8939, 1025.7739, 1025.6216, 1025.534, 1025.4138, 1025.3071, 1025.1984, 1025.0715, 1024.9052, 1024.7671, 1024.6786, 1024.4373, 1024.1082, 1024.0623, 1024.0359, 1023.99347, 1023.9526, 1023.9227, 1023.89886, 1023.8801, NaN, NaN, 1029.2588, 1029.2329, 1029.1969, 1029.1454, 1029.0953, 1029.0427, 1028.9924, 1028.9395, 1028.8905, 1028.8391, 1028.7927, 1028.7472, 1028.6951, 1028.6427, 1028.5869, 1028.5415, 1028.4946, 1028.4375, 1028.3792, 1028.3124, 1028.2579, 1028.208, 1028.1602, 1028.117, 1028.0752, 1028.0359, 1027.9911, 1027.9401, 1027.8906, 1027.845, 1027.7961, 1027.7482, 1027.6921, 1027.6367, 1027.5856, 1027.5411, 1027.4883, 1027.4324, 1027.382, 1027.3253, 1027.2618, 1027.2101, 1027.1383, 1027.0588, 1026.991, 1026.9292, 1026.8591, 1026.7639, 1026.6654, 1026.5774, 1026.4755, 1026.3185, 1026.1395, 1025.9607, 1025.7816, 1025.6311, 1025.507, 1025.3634, 1025.2341, 1025.104, 1024.9739, 1024.837, 1024.639, 1024.3905, 1024.2747, 1024.158, 1024.0446, 1023.98395, 1023.962, 1023.9418, 1023.92316, 1023.905, 1023.8837, 1023.8673, NaN, NaN, 1029.244, 1029.2166, 1029.181, 1029.1311, 1029.0817, 1029.0309, 1028.9774, 1028.933, 1028.8839, 1028.8331, 1028.7852, 1028.7429, 1028.6941, 1028.6528, 1028.6039, 1028.559, 1028.5063, 1028.4595, 1028.4088, 1028.3513, 1028.297, 1028.2412, 1028.1858, 1028.1318, 1028.0798, 1028.0352, 1027.9863, 1027.9425, 1027.8945, 1027.8441, 1027.7914, 1027.7401, 1027.6876, 1027.6338, 1027.5757, 1027.5297, 1027.4714, 1027.4056, 1027.3444, 1027.2776, 1027.21, 1027.1311, 1027.0345, 1026.9327, 1026.8247, 1026.7308, 1026.6304, 1026.5171, 1026.4219, 1026.262, 1026.145, 1025.981, 1025.8312, 1025.6732, 1025.5581, 1025.433, 1025.3245, 1025.2135, 1025.1393, 1025.0453, 1024.9391, 1024.7887, 1024.6124, 1024.4751, 1024.1409, 1024.0905, 1024.0664, 1024.0422, 1024.0157, 1023.98846, 1023.95667, 1023.93384, NaN, NaN, 1029.2681, 1029.2391, 1029.2042, 1029.1526, 1029.0942, 1029.0375, 1028.9823, 1028.9272, 1028.8724, 1028.8123, 1028.7576, 1028.7085, 1028.6631, 1028.6165, 1028.566, 1028.5205, 1028.4691, 1028.4148, 1028.3611, 1028.3013, 1028.2463, 1028.1918, 1028.1396, 1028.0848, 1028.0312, 1027.9794, 1027.9313, 1027.8762, 1027.8257, 1027.7769, 1027.713, 1027.6569, 1027.5997, 1027.5431, 1027.4829, 1027.4209, 1027.3586, 1027.2964, 1027.2261, 1027.1517, 1027.0775, 1026.9956, 1026.8832, 1026.7863, 1026.6748, 1026.593, 1026.4797, 1026.4053, 1026.2789, 1026.189, 1026.0706, 1025.9172, 1025.755, 1025.6385, 1025.5095, 1025.3873, 1025.2369, 1025.061, 1024.9219, 1024.802, 1024.6858, 1024.5387, 1024.3042, 1024.0287, 1023.9963, 1023.9732, 1023.94806, 1023.9203, 1023.8928, 1023.8743, NaN, NaN, 1029.2706, 1029.2432, 1029.2091, 1029.1536, 1029.1046, 1029.0594, 1029.0125, 1028.963, 1028.9042, 1028.8508, 1028.7998, 1028.7498, 1028.7028, 1028.6543, 1028.612, 1028.5707, 1028.5151, 1028.4666, 1028.4125, 1028.363, 1028.3121, 1028.2618, 1028.2107, 1028.1565, 1028.0986, 1028.0454, 1027.9908, 1027.9364, 1027.8707, 1027.8066, 1027.7473, 1027.6884, 1027.634, 1027.5664, 1027.4993, 1027.4348, 1027.3812, 1027.3263, 1027.2606, 1027.2008, 1027.1344, 1027.0532, 1026.9756, 1026.898, 1026.8152, 1026.7158, 1026.6184, 1026.4949, 1026.3552, 1026.2087, 1026.0665, 1025.9017, 1025.7456, 1025.5896, 1025.4254, 1025.3092, 1025.1414, 1025.019, 1024.8868, 1024.8032, 1024.5555, 1024.3153, 1024.0353, 1023.99207, 1023.9675, 1023.9454, 1023.91516, 1023.8955, 1023.8726, 1023.85864, NaN, NaN, 1029.2451, 1029.2118, 1029.1686, 1029.1157, 1029.0623, 1029.0073, 1028.954, 1028.8945, 1028.8397, 1028.7877, 1028.736, 1028.6885, 1028.6404, 1028.5957, 1028.554, 1028.5065, 1028.456, 1028.4095, 1028.355, 1028.3046, 1028.2568, 1028.208, 1028.1624, 1028.1156, 1028.0665, 1028.015, 1027.9667, 1027.912, 1027.8594, 1027.812, 1027.7546, 1027.7013, 1027.6455, 1027.594, 1027.5438, 1027.4968, 1027.4363, 1027.3629, 1027.301, 1027.2444, 1027.1882, 1027.1239, 1027.053, 1026.9866, 1026.9174, 1026.8582, 1026.7845, 1026.6727, 1026.5614, 1026.4502, 1026.2983, 1026.1968, 1026.0682, 1025.9128, 1025.7792, 1025.6552, 1025.4899, 1025.3605, 1025.2516, 1025.1097, 1025.036, 1024.9194, 1024.8276, 1024.6493, 1024.2408, 1024.0154, 1023.9957, 1023.97253, 1023.9504, 1023.9324, 1023.91016, 1023.8893, 1023.8683, NaN, NaN, 1029.2676, 1029.2416, 1029.2054, 1029.1523, 1029.1022, 1029.0513, 1029.0039, 1028.9503, 1028.8951, 1028.843, 1028.7819, 1028.7268, 1028.6726, 1028.6171, 1028.5663, 1028.5193, 1028.4735, 1028.4193, 1028.3624, 1028.3046, 1028.2546, 1028.2035, 1028.15, 1028.0991, 1028.049, 1028.001, 1027.9467, 1027.8893, 1027.832, 1027.776, 1027.7263, 1027.6774, 1027.624, 1027.5709, 1027.5087, 1027.4509, 1027.3993, 1027.3389, 1027.269, 1027.1879, 1027.116, 1027.0343, 1026.9645, 1026.8876, 1026.8108, 1026.7249, 1026.6171, 1026.4756, 1026.313, 1026.1687, 1026.0286, 1025.8671, 1025.6742, 1025.5154, 1025.4165, 1025.3646, 1025.2563, 1025.1221, 1024.9944, 1024.9202, 1024.748, 1024.5786, 1024.2931, 1024.1007, 1023.9852, 1023.9596, 1023.93414, 1023.9122, 1023.89294, 1023.8734, 1023.8535, NaN, NaN, 1029.2439, 1029.2145, 1029.1812, 1029.1329, 1029.0808, 1029.0306, 1028.982, 1028.9261, 1028.8759, 1028.8223, 1028.7699, 1028.7151, 1028.6646, 1028.6172, 1028.5659, 1028.5126, 1028.4628, 1028.4077, 1028.3594, 1028.3134, 1028.262, 1028.2083, 1028.1538, 1028.102, 1028.0519, 1027.9956, 1027.9421, 1027.8928, 1027.8403, 1027.7842, 1027.7239, 1027.6672, 1027.6147, 1027.5571, 1027.5004, 1027.447, 1027.3951, 1027.3268, 1027.2515, 1027.1628, 1027.0731, 1026.968, 1026.8663, 1026.7926, 1026.7083, 1026.5824, 1026.452, 1026.3141, 1026.168, 1026.0593, 1025.9185, 1025.798, 1025.6398, 1025.506, 1025.3867, 1025.2705, 1025.1416, 1025.0276, 1024.8243, 1024.5962, 1024.3114, 1024.0494, 1024.0061, 1023.98663, 1023.9618, 1023.9375, 1023.9152, 1023.891, 1023.8647, 1023.8409, 1023.83136, NaN, NaN, 1029.261, 1029.2338, 1029.1958, 1029.144, 1029.0994, 1029.0511, 1029.0015, 1028.9521, 1028.9042, 1028.8607, 1028.8086, 1028.7595, 1028.7081, 1028.655, 1028.6022, 1028.5533, 1028.5049, 1028.4619, 1028.4111, 1028.3531, 1028.3018, 1028.2524, 1028.2017, 1028.1488, 1028.0918, 1028.0358, 1027.9858, 1027.9376, 1027.8889, 1027.839, 1027.7858, 1027.7272, 1027.6755, 1027.6229, 1027.5686, 1027.5175, 1027.4608, 1027.4088, 1027.3567, 1027.2913, 1027.2169, 1027.1332, 1027.0483, 1026.9689, 1026.889, 1026.8036, 1026.719, 1026.5934, 1026.467, 1026.3599, 1026.2557, 1026.0989, 1025.9237, 1025.7675, 1025.56, 1025.4752, 1025.3318, 1025.2158, 1025.1273, 1025.0161, 1024.8782, 1024.7423, 1024.5187, 1024.1156, 1024.0138, 1023.9936, 1023.9734, 1023.949, 1023.927, 1023.9023, 1023.8836, NaN, NaN, 1029.2551, 1029.2278, 1029.1898, 1029.1394, 1029.0853, 1029.0345, 1028.9838, 1028.9348, 1028.8833, 1028.8333, 1028.7811, 1028.7297, 1028.6748, 1028.6233, 1028.5692, 1028.518, 1028.4698, 1028.4182, 1028.3707, 1028.32, 1028.2623, 1028.2112, 1028.1593, 1028.1108, 1028.0579, 1028.0093, 1027.9554, 1027.901, 1027.8534, 1027.7996, 1027.7411, 1027.6847, 1027.6326, 1027.5754, 1027.5259, 1027.4703, 1027.4111, 1027.3539, 1027.285, 1027.2227, 1027.1527, 1027.0745, 1027.0018, 1026.9294, 1026.8086, 1026.6969, 1026.571, 1026.4741, 1026.3516, 1026.2126, 1026.0558, 1025.959, 1025.8276, 1025.6873, 1025.5585, 1025.4442, 1025.3353, 1025.2842, 1025.1952, 1025.1118, 1024.9789, 1024.7863, 1024.629, 1024.3434, 1024.0056, 1023.9877, 1023.97253, 1023.9509, 1023.9271, 1023.9094, 1023.8906, 1023.871, 1023.8568, NaN, NaN, 1029.2307, 1029.2042, 1029.1672, 1029.1211, 1029.0729, 1029.0256, 1028.9772, 1028.9269, 1028.875, 1028.819, 1028.7711, 1028.721, 1028.6663, 1028.6067, 1028.5509, 1028.5037, 1028.4541, 1028.3995, 1028.3478, 1028.2919, 1028.2255, 1028.1677, 1028.1144, 1028.0605, 1027.9985, 1027.9495, 1027.899, 1027.8447, 1027.7839, 1027.7277, 1027.6747, 1027.623, 1027.5789, 1027.5269, 1027.4691, 1027.4147, 1027.357, 1027.3033, 1027.2246, 1027.167, 1027.098, 1027.0299, 1026.9268, 1026.8253, 1026.714, 1026.5972, 1026.4978, 1026.4208, 1026.3275, 1026.1808, 1026.0139, 1025.8982, 1025.776, 1025.6318, 1025.4503, 1025.3357, 1025.2502, 1025.1334, 1025.0021, 1024.8239, 1024.6359, 1024.2769, 1024.0277, 1024.0095, 1023.9893, 1023.96906, 1023.95135, 1023.92505, 1023.89844, 1023.8849, NaN, NaN, 1029.2273, 1029.1978, 1029.1619, 1029.1075, 1029.0541, 1029.0034, 1028.9519, 1028.9004, 1028.852, 1028.8, 1028.744, 1028.6906, 1028.6398, 1028.5814, 1028.5332, 1028.4846, 1028.4321, 1028.3811, 1028.3254, 1028.2731, 1028.22, 1028.1663, 1028.1238, 1028.0731, 1028.0117, 1027.9587, 1027.9045, 1027.8425, 1027.7863, 1027.7395, 1027.6926, 1027.639, 1027.5815, 1027.5253, 1027.4731, 1027.4111, 1027.3522, 1027.2937, 1027.2284, 1027.1594, 1027.0929, 1027.0251, 1026.9423, 1026.8502, 1026.7411, 1026.6317, 1026.5288, 1026.4393, 1026.2725, 1026.0923, 1025.9291, 1025.7986, 1025.6041, 1025.4319, 1025.3408, 1025.2446, 1025.1295, 1025.0144, 1024.8921, 1024.7554, 1024.5071, 1024.2739, 1024.0251, 1024.002, 1023.9782, 1023.95483, 1023.9299, 1023.9071, 1023.8886, 1023.8658, NaN, NaN, 1029.2173, 1029.1886, 1029.1537, 1029.1115, 1029.0623, 1029.011, 1028.961, 1028.9141, 1028.8643, 1028.8129, 1028.7621, 1028.714, 1028.6661, 1028.6187, 1028.5702, 1028.527, 1028.4824, 1028.4374, 1028.3905, 1028.3372, 1028.288, 1028.2393, 1028.1913, 1028.1412, 1028.0931, 1028.0417, 1027.9924, 1027.9421, 1027.8842, 1027.8254, 1027.7648, 1027.7089, 1027.6519, 1027.5991, 1027.5452, 1027.4927, 1027.438, 1027.3871, 1027.3378, 1027.2863, 1027.2203, 1027.156, 1027.0598, 1026.9773, 1026.9014, 1026.8094, 1026.691, 1026.6091, 1026.4884, 1026.3645, 1026.2012, 1026.0372, 1025.8342, 1025.7106, 1025.5704, 1025.4619, 1025.3496, 1025.2261, 1025.1215, 1025.0149, 1024.89, 1024.7721, 1024.5607, 1024.2925, 1024.0789, 1024.0536, 1024.0295, 1024.0112, 1023.98755, 1023.9646, 1023.9462, 1023.9249, 1023.9058, 1023.88446, NaN, NaN, 1029.232, 1029.2063, 1029.1688, 1029.1199, 1029.0736, 1029.0256, 1028.9727, 1028.9272, 1028.8771, 1028.8247, 1028.7732, 1028.7246, 1028.6743, 1028.6284, 1028.5831, 1028.5342, 1028.4835, 1028.4368, 1028.3881, 1028.3364, 1028.2876, 1028.2351, 1028.1768, 1028.1198, 1028.0594, 1028.0106, 1027.9514, 1027.9008, 1027.844, 1027.7947, 1027.7433, 1027.694, 1027.6438, 1027.5847, 1027.5292, 1027.4747, 1027.4202, 1027.3533, 1027.2968, 1027.234, 1027.168, 1027.0997, 1027.0338, 1026.9679, 1026.8611, 1026.7611, 1026.6823, 1026.5831, 1026.481, 1026.2876, 1026.1827, 1026.0415, 1025.9297, 1025.7759, 1025.6289, 1025.4468, 1025.3127, 1025.1561, 1025.0547, 1024.8827, 1024.6271, 1024.2491, 1024.0647, 1024.0403, 1024.017, 1023.9905, 1023.96545, 1023.93677, 1023.9141, 1023.89276, 1023.86597, NaN, NaN, 1029.2308, 1029.2051, 1029.1697, 1029.1227, 1029.0708, 1029.0201, 1028.9684, 1028.9178, 1028.8688, 1028.8228, 1028.7727, 1028.72, 1028.6685, 1028.6141, 1028.5669, 1028.5132, 1028.4657, 1028.4211, 1028.369, 1028.3169, 1028.2678, 1028.2068, 1028.1571, 1028.1068, 1028.0553, 1028.0037, 1027.945, 1027.8873, 1027.8285, 1027.7776, 1027.7195, 1027.6631, 1027.6057, 1027.5435, 1027.478, 1027.4192, 1027.3644, 1027.2893, 1027.2126, 1027.1555, 1027.085, 1027.0269, 1026.9501, 1026.8629, 1026.7721, 1026.7054, 1026.6255, 1026.5168, 1026.417, 1026.3297, 1026.2471, 1026.0842, 1025.9613, 1025.799, 1025.6571, 1025.5221, 1025.3654, 1025.1924, 1025.0604, 1024.8757, 1024.66, 1024.1348, 1024.0604, 1024.0388, 1024.0168, 1023.9988, 1023.97186, 1023.943, 1023.9318, 1023.9153, 1023.89795, 1023.8701, NaN, NaN, 1029.2201, 1029.195, 1029.156, 1029.1086, 1029.0605, 1029.0076, 1028.9585, 1028.9088, 1028.8574, 1028.8087, 1028.7632, 1028.7142, 1028.6659, 1028.6161, 1028.5615, 1028.5096, 1028.4598, 1028.4127, 1028.3634, 1028.3167, 1028.2606, 1028.2019, 1028.1523, 1028.1031, 1028.0531, 1027.9988, 1027.944, 1027.8967, 1027.8398, 1027.7854, 1027.7357, 1027.6754, 1027.6201, 1027.5746, 1027.524, 1027.4696, 1027.414, 1027.3516, 1027.2878, 1027.2262, 1027.1609, 1027.0964, 1027.0382, 1026.9722, 1026.8778, 1026.7708, 1026.6808, 1026.5863, 1026.4667, 1026.3435, 1026.2085, 1026.0995, 1025.9435, 1025.8195, 1025.736, 1025.5952, 1025.481, 1025.3485, 1025.2377, 1025.1184, 1024.9933, 1024.8903, 1024.7375, 1024.5204, 1024.0267, 1024.0068, 1023.98285, 1023.958, 1023.93634, 1023.9144, 1023.88513, 1023.86066, NaN, NaN, 1029.2244, 1029.1979, 1029.1604, 1029.1128, 1029.0712, 1029.0194, 1028.97, 1028.921, 1028.866, 1028.8167, 1028.767, 1028.7126, 1028.6614, 1028.6122, 1028.558, 1028.4998, 1028.4435, 1028.3943, 1028.3468, 1028.2986, 1028.2488, 1028.2007, 1028.1487, 1028.09, 1028.0319, 1027.9792, 1027.9279, 1027.88, 1027.8287, 1027.771, 1027.7135, 1027.6531, 1027.5924, 1027.5433, 1027.4846, 1027.4279, 1027.3682, 1027.308, 1027.2344, 1027.1483, 1027.0731, 1027.002, 1026.9304, 1026.8462, 1026.7607, 1026.6534, 1026.5222, 1026.4412, 1026.33, 1026.144, 1025.9329, 1025.7885, 1025.6918, 1025.5116, 1025.4137, 1025.2932, 1025.1871, 1025.06, 1024.9526, 1024.808, 1024.6246, 1024.1989, 1024.0232, 1024.0032, 1023.98267, 1023.95856, 1023.93463, 1023.9134, 1023.89264, 1023.87317, 1023.8588, NaN, NaN, 1029.2219, 1029.1941, 1029.1556, 1029.11, 1029.0607, 1029.0161, 1028.9689, 1028.9227, 1028.8723, 1028.8278, 1028.7809, 1028.7308, 1028.6782, 1028.6279, 1028.5769, 1028.528, 1028.4788, 1028.4269, 1028.3789, 1028.3281, 1028.2771, 1028.2266, 1028.1782, 1028.1292, 1028.0747, 1028.0208, 1027.9645, 1027.9161, 1027.8693, 1027.8156, 1027.7646, 1027.7122, 1027.6567, 1027.6139, 1027.5514, 1027.5012, 1027.4424, 1027.3833, 1027.3177, 1027.2577, 1027.1877, 1027.1195, 1027.0421, 1026.959, 1026.8824, 1026.7891, 1026.6973, 1026.5792, 1026.4591, 1026.3654, 1026.1677, 1026.0217, 1025.8827, 1025.7599, 1025.7079, 1025.5997, 1025.483, 1025.35, 1025.2296, 1025.1094, 1024.9111, 1024.7555, 1024.47, 1024.0236, 1023.99994, 1023.98157, 1023.96814, 1023.953, 1023.9316, 1023.9132, 1023.88965, 1023.8674, 1023.8452, NaN, NaN, 1029.2327, 1029.2026, 1029.1643, 1029.1145, 1029.0594, 1029.0063, 1028.9517, 1028.9047, 1028.8501, 1028.7991, 1028.7506, 1028.6971, 1028.6406, 1028.5898, 1028.5403, 1028.4889, 1028.4337, 1028.38, 1028.3279, 1028.2698, 1028.2153, 1028.1558, 1028.0972, 1028.0453, 1027.9951, 1027.937, 1027.8802, 1027.8264, 1027.767, 1027.7148, 1027.6584, 1027.602, 1027.5417, 1027.4863, 1027.4226, 1027.3676, 1027.303, 1027.2317, 1027.1661, 1027.1069, 1027.0393, 1026.95, 1026.8629, 1026.7672, 1026.6992, 1026.6173, 1026.4392, 1026.2896, 1026.1722, 1026.0461, 1025.8616, 1025.7208, 1025.6155, 1025.491, 1025.402, 1025.2528, 1025.1058, 1024.9878, 1024.9067, 1024.7441, 1024.3585, 1024.0063, 1023.98505, 1023.9632, 1023.94476, 1023.92944, 1023.9138, 1023.8939, 1023.8684, 1023.8517, NaN, NaN, 1029.2368, 1029.2112, 1029.1729, 1029.1241, 1029.0819, 1029.0403, 1028.9923, 1028.9465, 1028.8966, 1028.856, 1028.8073, 1028.7552, 1028.7008, 1028.6492, 1028.5964, 1028.5485, 1028.497, 1028.443, 1028.3867, 1028.338, 1028.2872, 1028.2346, 1028.181, 1028.1235, 1028.0707, 1028.021, 1027.9648, 1027.9082, 1027.8544, 1027.806, 1027.753, 1027.7003, 1027.6444, 1027.5886, 1027.5286, 1027.4745, 1027.4197, 1027.3624, 1027.3021, 1027.2423, 1027.1774, 1027.1067, 1027.0422, 1026.9589, 1026.8582, 1026.7704, 1026.6838, 1026.6049, 1026.5242, 1026.4213, 1026.2792, 1026.0677, 1025.8555, 1025.7018, 1025.5708, 1025.4065, 1025.263, 1025.1716, 1025.0974, 1024.9911, 1024.8497, 1024.6458, 1024.136, 1024.0306, 1024.0134, 1023.99713, 1023.97943, 1023.9599, 1023.9368, 1023.9137, 1023.89026, 1023.86676, 1023.854, NaN, NaN, 1029.2153, 1029.1868, 1029.1525, 1029.104, 1029.0599, 1029.011, 1028.9597, 1028.9175, 1028.8662, 1028.8206, 1028.7748, 1028.7214, 1028.6785, 1028.6261, 1028.5767, 1028.53, 1028.4801, 1028.4312, 1028.3767, 1028.3254, 1028.2728, 1028.2183, 1028.165, 1028.1066, 1028.0547, 1028.0066, 1027.9545, 1027.9043, 1027.8561, 1027.8035, 1027.7521, 1027.6973, 1027.6373, 1027.5896, 1027.5371, 1027.4786, 1027.4271, 1027.3716, 1027.3086, 1027.2467, 1027.1884, 1027.1117, 1027.0311, 1026.9521, 1026.8691, 1026.7915, 1026.7035, 1026.6265, 1026.5254, 1026.4069, 1026.2279, 1026.069, 1025.9198, 1025.7759, 1025.6288, 1025.4987, 1025.3329, 1025.2434, 1025.1464, 1025.0143, 1024.8491, 1024.7438, 1024.6672, 1024.2998, 1024.0292, 1024.0117, 1023.98785, 1023.9658, 1023.94574, 1023.9221, 1023.90186, 1023.8791, 1023.86053, NaN, NaN, 1029.2196, 1029.1942, 1029.1525, 1029.1077, 1029.0587, 1029.0095, 1028.9563, 1028.9108, 1028.8586, 1028.8094, 1028.7583, 1028.7074, 1028.6587, 1028.6102, 1028.5631, 1028.5088, 1028.4604, 1028.4156, 1028.3666, 1028.3116, 1028.261, 1028.2104, 1028.1552, 1028.1086, 1028.0564, 1028.0077, 1027.9623, 1027.9117, 1027.8647, 1027.8102, 1027.7548, 1027.7078, 1027.6592, 1027.6069, 1027.5596, 1027.5092, 1027.4424, 1027.3889, 1027.3331, 1027.2607, 1027.1796, 1027.1072, 1027.0343, 1026.9451, 1026.8503, 1026.7649, 1026.6646, 1026.5518, 1026.4424, 1026.3337, 1026.2151, 1026.0947, 1025.9491, 1025.8013, 1025.6787, 1025.5781, 1025.4591, 1025.3274, 1025.2225, 1025.1127, 1025.0076, 1024.8882, 1024.7716, 1024.64, 1024.4888, 1024.131, 1024.0245, 1023.984, 1023.9609, 1023.93805, 1023.9171, 1023.89355, 1023.8653, 1023.8425, NaN, NaN, 1029.2084, 1029.18, 1029.1411, 1029.0874, 1029.0309, 1028.9757, 1028.92, 1028.8634, 1028.8092, 1028.7545, 1028.6995, 1028.6477, 1028.5956, 1028.5375, 1028.4906, 1028.4419, 1028.3889, 1028.3385, 1028.2869, 1028.2356, 1028.1765, 1028.121, 1028.0717, 1028.0126, 1027.9563, 1027.9025, 1027.846, 1027.793, 1027.739, 1027.6871, 1027.6299, 1027.5784, 1027.5236, 1027.4674, 1027.4072, 1027.3472, 1027.2834, 1027.2269, 1027.1597, 1027.0852, 1027.0212, 1026.948, 1026.858, 1026.7638, 1026.6539, 1026.5548, 1026.4696, 1026.4015, 1026.3058, 1026.1663, 1026.0474, 1025.8818, 1025.7349, 1025.5942, 1025.51, 1025.3508, 1025.2432, 1025.1813, 1025.0929, 1025.028, 1024.9384, 1024.8081, 1024.5626, 1024.1611, 1024.0001, 1023.9765, 1023.951, 1023.9289, 1023.90295, 1023.8791, 1023.8494, NaN, NaN, 1029.2322, 1029.2067, 1029.1691, 1029.1243, 1029.0702, 1029.0199, 1028.9753, 1028.9274, 1028.88, 1028.8385, 1028.7859, 1028.7338, 1028.6858, 1028.6364, 1028.588, 1028.5391, 1028.4844, 1028.4332, 1028.386, 1028.3376, 1028.2854, 1028.231, 1028.1802, 1028.1266, 1028.0841, 1028.0433, 1028.0024, 1027.9625, 1027.9229, 1027.8871, 1027.8457, 1027.809, 1027.7751, 1027.7375, 1027.703, 1027.6636, 1027.6215, 1027.5731, 1027.5211, 1027.4612, 1027.412, 1027.3674, 1027.3206, 1027.2635, 1027.2104, 1027.1594, 1027.0996, 1027.047, 1026.9911, 1026.9247, 1026.8497, 1026.7709, 1026.6858, 1026.5846, 1026.4525, 1026.3453, 1026.246, 1026.1118, 1025.9402, 1025.8123, 1025.709, 1025.5825, 1025.4338, 1025.3275, 1025.2074, 1025.1003, 1024.9694, 1024.7485, 1024.4412, 1024.1251, 1024.0538, 1024.0276, 1024.0012, 1023.97766, 1023.9537, 1023.93, 1023.9036, 1023.8742, 1023.8538, NaN, NaN, 1029.2468, 1029.2196, 1029.1815, 1029.1277, 1029.0754, 1029.0259, 1028.9752, 1028.929, 1028.878, 1028.826, 1028.7731, 1028.7179, 1028.669, 1028.6184, 1028.5657, 1028.5123, 1028.4624, 1028.4099, 1028.36, 1028.3165, 1028.27, 1028.2205, 1028.1742, 1028.1235, 1028.0737, 1028.02, 1027.9717, 1027.9194, 1027.8691, 1027.8148, 1027.7681, 1027.7094, 1027.6548, 1027.6029, 1027.556, 1027.5005, 1027.4375, 1027.3732, 1027.3094, 1027.2487, 1027.188, 1027.1224, 1027.0538, 1026.992, 1026.9208, 1026.837, 1026.7524, 1026.6436, 1026.5133, 1026.3755, 1026.2344, 1026.0724, 1025.8888, 1025.7157, 1025.5806, 1025.4285, 1025.2838, 1025.1525, 1025.0636, 1024.9863, 1024.8013, 1024.5521, 1024.2155, 1024.0718, 1024.0474, 1024.0215, 1023.99225, 1023.95685, 1023.9272, 1023.898, 1023.8764, NaN, NaN, 1029.2155, 1029.1849, 1029.1494, 1029.0973, 1029.044, 1028.9908, 1028.9391, 1028.8917, 1028.8359, 1028.7843, 1028.7341, 1028.6906, 1028.6443, 1028.598, 1028.5543, 1028.5045, 1028.4543, 1028.4012, 1028.3441, 1028.2892, 1028.241, 1028.1946, 1028.1416, 1028.0944, 1028.0486, 1027.9994, 1027.9489, 1027.8992, 1027.8507, 1027.7947, 1027.7395, 1027.6871, 1027.6366, 1027.5779, 1027.529, 1027.4767, 1027.42, 1027.3611, 1027.2964, 1027.2341, 1027.1573, 1027.094, 1027.0232, 1026.952, 1026.8735, 1026.7856, 1026.7046, 1026.5958, 1026.4788, 1026.3655, 1026.2053, 1026.0453, 1025.8661, 1025.7067, 1025.597, 1025.476, 1025.4133, 1025.3, 1025.2272, 1025.1384, 1025.0273, 1024.887, 1024.7374, 1024.5613, 1024.3945, 1024.0925, 1024.0704, 1024.0463, 1024.0238, 1023.999, 1023.96674, 1023.92914, 1023.901, 1023.88715, NaN, NaN, 1029.2151, 1029.1808, 1029.1465, 1029.0946, 1029.0441, 1028.9894, 1028.9336, 1028.8773, 1028.8265, 1028.7787, 1028.7308, 1028.6812, 1028.6339, 1028.5817, 1028.5354, 1028.4885, 1028.4377, 1028.3856, 1028.3352, 1028.2839, 1028.2336, 1028.1816, 1028.132, 1028.0785, 1028.034, 1027.9829, 1027.9287, 1027.877, 1027.8203, 1027.7595, 1027.7076, 1027.6516, 1027.5974, 1027.5385, 1027.485, 1027.4346, 1027.368, 1027.3024, 1027.2383, 1027.167, 1027.1036, 1027.035, 1026.96, 1026.8806, 1026.8241, 1026.7377, 1026.6603, 1026.5754, 1026.4491, 1026.3015, 1026.1525, 1026.0371, 1025.883, 1025.7969, 1025.6752, 1025.568, 1025.4487, 1025.351, 1025.2346, 1025.1356, 1025.0208, 1024.8773, 1024.7041, 1024.5011, 1024.3221, 1024.0948, 1024.0406, 1024.0142, 1023.99023, 1023.9656, 1023.9385, 1023.91455, 1023.8978, NaN, NaN, 1029.2479, 1029.2177, 1029.177, 1029.1255, 1029.0767, 1029.0289, 1028.9756, 1028.9259, 1028.8721, 1028.8147, 1028.7648, 1028.7188, 1028.6658, 1028.6151, 1028.5663, 1028.5214, 1028.4755, 1028.4257, 1028.375, 1028.3236, 1028.2725, 1028.2241, 1028.1724, 1028.1285, 1028.0793, 1028.0262, 1027.9714, 1027.9154, 1027.8552, 1027.805, 1027.7509, 1027.6952, 1027.6404, 1027.5908, 1027.5392, 1027.4828, 1027.4197, 1027.3617, 1027.2858, 1027.2208, 1027.1581, 1027.0953, 1027.0264, 1026.9614, 1026.8947, 1026.8219, 1026.7446, 1026.6742, 1026.5706, 1026.4551, 1026.3358, 1026.2, 1026.0697, 1025.9197, 1025.7811, 1025.6339, 1025.4893, 1025.3522, 1025.2329, 1025.0953, 1025.014, 1024.8959, 1024.7554, 1024.5149, 1024.2708, 1024.1141, 1024.07, 1024.0487, 1024.0271, 1024.0055, 1023.98346, 1023.95856, 1023.93616, NaN, NaN, 1029.2053, 1029.1798, 1029.1478, 1029.105, 1029.0636, 1029.0173, 1028.9692, 1028.926, 1028.8794, 1028.8403, 1028.7903, 1028.7466, 1028.7034, 1028.6573, 1028.6113, 1028.5669, 1028.5225, 1028.476, 1028.4264, 1028.3755, 1028.3263, 1028.2767, 1028.2208, 1028.1675, 1028.1163, 1028.0723, 1028.0309, 1027.9839, 1027.9359, 1027.8877, 1027.839, 1027.7875, 1027.7386, 1027.6937, 1027.6407, 1027.5895, 1027.5406, 1027.4923, 1027.4324, 1027.3876, 1027.3193, 1027.246, 1027.1876, 1027.1134, 1027.0486, 1026.9775, 1026.9093, 1026.8417, 1026.7717, 1026.6918, 1026.6302, 1026.5446, 1026.4296, 1026.3373, 1026.2277, 1026.0934, 1025.9049, 1025.7625, 1025.6119, 1025.4519, 1025.3365, 1025.2151, 1025.1282, 1024.9854, 1024.7777, 1024.429, 1024.2659, 1024.1487, 1024.1046, 1024.082, 1024.06, 1024.0369, 1024.0175, 1023.9911, 1023.9658, 1023.9446, 1023.9297, NaN, NaN, 1029.2201, 1029.1938, 1029.1613, 1029.1151, 1029.0706, 1029.0278, 1028.9827, 1028.9373, 1028.889, 1028.8418, 1028.795, 1028.7513, 1028.7045, 1028.6567, 1028.6074, 1028.5625, 1028.5114, 1028.4646, 1028.42, 1028.3733, 1028.321, 1028.2727, 1028.2195, 1028.1692, 1028.1179, 1028.0757, 1028.0344, 1027.9875, 1027.9415, 1027.896, 1027.8438, 1027.7944, 1027.7456, 1027.6958, 1027.6439, 1027.586, 1027.5367, 1027.4768, 1027.4132, 1027.3604, 1027.292, 1027.2365, 1027.1533, 1027.0742, 1026.9944, 1026.9302, 1026.8646, 1026.7771, 1026.6807, 1026.5844, 1026.4849, 1026.3525, 1026.1885, 1026.0822, 1025.9364, 1025.7643, 1025.6262, 1025.4885, 1025.3549, 1025.2434, 1025.1147, 1024.9382, 1024.6967, 1024.4452, 1024.2758, 1024.1915, 1024.0797, 1024.0576, 1024.0343, 1024.0116, 1023.9895, 1023.96783, 1023.94324, 1023.9223, NaN, NaN, 1029.1968, 1029.1697, 1029.1335, 1029.0868, 1029.0425, 1028.9951, 1028.946, 1028.8986, 1028.85, 1028.8037, 1028.7554, 1028.7068, 1028.653, 1028.6074, 1028.5642, 1028.5155, 1028.4628, 1028.4083, 1028.3545, 1028.3042, 1028.2499, 1028.2039, 1028.1552, 1028.1011, 1028.0466, 1027.9908, 1027.9412, 1027.8911, 1027.8424, 1027.7903, 1027.7365, 1027.6868, 1027.6301, 1027.5739, 1027.5267, 1027.4755, 1027.4185, 1027.3613, 1027.2965, 1027.2415, 1027.161, 1027.0801, 1027.0073, 1026.9229, 1026.8567, 1026.772, 1026.6853, 1026.5807, 1026.471, 1026.3754, 1026.2186, 1026.0948, 1025.9993, 1025.8741, 1025.7474, 1025.606, 1025.4838, 1025.337, 1025.2003, 1025.1027, 1024.9916, 1024.8774, 1024.7296, 1024.565, 1024.307, 1024.1517, 1024.063, 1024.0432, 1024.021, 1024.0, 1023.9769, 1023.9545, 1023.9307, 1023.90686, NaN, NaN, 1029.209, 1029.1808, 1029.1467, 1029.1017, 1029.0605, 1029.019, 1028.9746, 1028.9287, 1028.8849, 1028.8407, 1028.7971, 1028.7543, 1028.7053, 1028.661, 1028.6182, 1028.5734, 1028.5347, 1028.4851, 1028.4364, 1028.394, 1028.3453, 1028.3, 1028.2518, 1028.2053, 1028.1611, 1028.1111, 1028.0651, 1028.0214, 1027.9656, 1027.9144, 1027.8622, 1027.8098, 1027.7607, 1027.7115, 1027.6573, 1027.6063, 1027.5642, 1027.5096, 1027.4507, 1027.3966, 1027.3469, 1027.2815, 1027.2205, 1027.146, 1027.0757, 1026.9944, 1026.9215, 1026.857, 1026.7689, 1026.6808, 1026.558, 1026.3983, 1026.2848, 1026.2137, 1026.1005, 1025.9711, 1025.9188, 1025.7659, 1025.6051, 1025.4988, 1025.3658, 1025.2502, 1025.1315, 1025.0176, 1024.8761, 1024.7228, 1024.4196, 1024.2343, 1024.1157, 1024.0853, 1024.061, 1024.0359, 1024.0072, 1023.9795, 1023.9478, 1023.9144, 1023.88983, NaN, NaN, 1029.2162, 1029.1902, 1029.1567, 1029.1073, 1029.0541, 1029.0046, 1028.9576, 1028.9021, 1028.8512, 1028.8007, 1028.7501, 1028.6962, 1028.648, 1028.6045, 1028.5546, 1028.5033, 1028.449, 1028.4058, 1028.3575, 1028.3136, 1028.271, 1028.22, 1028.1713, 1028.1208, 1028.07, 1028.0243, 1027.9801, 1027.9252, 1027.8722, 1027.8223, 1027.7726, 1027.7211, 1027.6747, 1027.6224, 1027.5681, 1027.518, 1027.4586, 1027.3906, 1027.3317, 1027.2745, 1027.2174, 1027.1584, 1027.0752, 1026.9888, 1026.9105, 1026.8392, 1026.7664, 1026.6813, 1026.5704, 1026.4333, 1026.2839, 1026.132, 1026.0045, 1025.8618, 1025.7133, 1025.5725, 1025.4735, 1025.3566, 1025.2263, 1025.0825, 1024.9069, 1024.7751, 1024.3569, 1024.1948, 1024.106, 1024.0819, 1024.0625, 1024.0388, 1024.0194, 1023.99774, 1023.9712, 1023.9419, 1023.90234, 1023.881, NaN, NaN, 1029.2208, 1029.1919, 1029.1572, 1029.1058, 1029.0537, 1028.9993, 1028.9464, 1028.8969, 1028.8456, 1028.7936, 1028.749, 1028.6956, 1028.6482, 1028.592, 1028.5431, 1028.4924, 1028.4415, 1028.3926, 1028.3363, 1028.2887, 1028.2311, 1028.1766, 1028.1229, 1028.0681, 1028.0148, 1027.966, 1027.9119, 1027.8608, 1027.8075, 1027.7578, 1027.7102, 1027.6572, 1027.596, 1027.535, 1027.4789, 1027.4104, 1027.3473, 1027.2708, 1027.2017, 1027.1516, 1027.0868, 1027.0054, 1026.9231, 1026.8354, 1026.7695, 1026.6869, 1026.5762, 1026.4697, 1026.3616, 1026.1993, 1026.0181, 1025.8524, 1025.7189, 1025.6097, 1025.4933, 1025.3993, 1025.2297, 1025.0627, 1024.9105, 1024.7894, 1024.5665, 1024.2607, 1024.127, 1024.0615, 1024.0391, 1024.0148, 1023.99005, 1023.96295, 1023.93555, 1023.9122, 1023.8991, NaN, NaN, 1029.2064, 1029.1743, 1029.1383, 1029.088, 1029.0424, 1028.9955, 1028.9456, 1028.9004, 1028.852, 1028.8091, 1028.765, 1028.7223, 1028.6791, 1028.6346, 1028.5918, 1028.5437, 1028.5005, 1028.4487, 1028.3982, 1028.3479, 1028.3, 1028.2571, 1028.2053, 1028.156, 1028.1027, 1028.0626, 1028.0114, 1027.9617, 1027.9141, 1027.8685, 1027.8196, 1027.7654, 1027.7163, 1027.6697, 1027.6234, 1027.569, 1027.5143, 1027.4542, 1027.4, 1027.3463, 1027.2922, 1027.2312, 1027.1671, 1027.098, 1027.0244, 1026.9713, 1026.8934, 1026.8052, 1026.6982, 1026.592, 1026.5125, 1026.4346, 1026.302, 1026.1554, 1026.0392, 1025.8774, 1025.7778, 1025.6423, 1025.485, 1025.4216, 1025.3184, 1025.1761, 1025.052, 1024.8707, 1024.7256, 1024.396, 1024.1143, 1024.0718, 1024.051, 1024.025, 1024.002, 1023.9814, 1023.9572, 1023.9346, 1023.9168, NaN, NaN, 1029.2069, 1029.18, 1029.145, 1029.0975, 1029.0563, 1029.0117, 1028.9681, 1028.9216, 1028.874, 1028.8293, 1028.7793, 1028.7313, 1028.6816, 1028.6338, 1028.5905, 1028.5388, 1028.4918, 1028.4386, 1028.3828, 1028.3353, 1028.291, 1028.243, 1028.1931, 1028.1464, 1028.099, 1028.0422, 1027.9874, 1027.9369, 1027.886, 1027.8342, 1027.7836, 1027.7333, 1027.676, 1027.6295, 1027.5818, 1027.5336, 1027.4817, 1027.4336, 1027.3833, 1027.3323, 1027.2771, 1027.2039, 1027.1354, 1027.0619, 1026.9789, 1026.9038, 1026.8024, 1026.7017, 1026.603, 1026.4729, 1026.3754, 1026.2306, 1026.0695, 1025.9377, 1025.7937, 1025.6416, 1025.5077, 1025.4318, 1025.3221, 1025.229, 1025.1411, 1025.0007, 1024.9229, 1024.8134, 1024.6576, 1024.4443, 1024.1226, 1024.0347, 1024.0093, 1023.987, 1023.9613, 1023.93896, 1023.91986, 1023.89813, NaN}
    DOXY = 
      {NaN, 115.05980666088254, 113.07850013591418, 111.6825719100918, 110.5070220081778, 109.84324347745851, 109.40022898751432, 109.1419418994265, 109.36169187786409, 110.77929699628912, 111.75965292100236, 113.67695736676589, 115.87205917215722, 117.79566005282652, 120.01828530960017, 121.93641789349844, 124.20661000269233, 125.06299576346422, 126.10154449508404, 126.06916154742689, 125.60681919069803, 124.54411190629457, 123.2222665488057, 121.23882293370986, 118.60000789351204, 116.84561906810727, 114.31731983021426, 113.0002877582427, 112.78722245301438, 114.22865066111441, 115.10186380374611, 115.97869288875096, 116.63246013165438, 116.9548309645072, 117.50116503707716, 118.93174480286038, 122.02246541239292, 126.77690220278096, 130.53074353191826, 138.38717629782505, 149.65703428203872, 157.11649358189328, 166.04332171004748, 171.42309998243917, 176.71812673940215, 182.1135986834304, 186.72785911515857, 191.84829251856692, 196.8120648455679, 199.54073232564187, 202.415383375781, 204.19319862254926, 205.81568365686698, 208.28571980185356, 210.02280554143422, 212.70167817754654, 216.71531365429132, 218.65063484883288, 220.19091305694246, 221.28954023017886, 220.38882630706684, 222.7480915547292, 222.96332076479592, 221.44301990954696, 221.95631168855274, 227.32141282878695, 231.5040494781019, 235.13745941286902, 239.06010790486985, 242.3308658973293, 247.0179726340796, 251.15254274080382, 253.49970298360898, 255.7763814111332, 257.23467568142934, 258.03039352040906, 258.9075863670458, 259.26511903617285, 259.8435355515475, 260.1320926701702, NaN, NaN, 118.66530851566847, 115.7311189859348, 113.27276837036565, 111.94984257111682, 112.44883630591347, 113.62298096195467, 115.29413127891513, 116.1056956349858, 117.16898124491031, 117.89990171344441, 118.55877375348238, 119.29637477401661, 119.95877864526483, 120.7024945855073, 121.78173726880804, 123.47651536203519, 124.61175859949371, 125.61175273970146, 125.75709853868379, 123.3431228300398, 120.72238465623788, 118.37678283614365, 116.32501470861416, 114.63826771786363, 114.16597145575889, 114.05438971070471, 113.90320947377352, 113.34889583358559, 113.45968608312577, 116.24328651807201, 119.2200269804151, 122.26416273770008, 123.68963619837886, 125.37579467651672, 126.47009277655249, 127.49438099678677, 129.06806064372668, 130.45884602094756, 132.96113015448287, 134.95353110466434, 137.01014257219603, 142.37861385131225, 146.13440823182142, 154.52326758119898, 160.29238751358184, 165.29374082728046, 169.33331677910655, 171.83337041150153, 174.6332086724282, 178.69156937519108, 182.0163294782881, 186.23321239613685, 190.0913235470776, 193.86304253568332, 198.50484047639088, 201.80102649005033, 204.916588848531, 209.15729696568104, 211.6852675391817, 214.33721444902753, 217.27962023468552, 216.2597636005569, 216.5136090679196, 218.99292821161742, 223.12205349922593, 230.71834342142225, 234.56013985225508, 238.49527967759394, 243.07856132867354, 246.41823904796112, 249.36371882567127, 251.6407874478767, 253.47503073299288, 254.94105540431045, 256.2545410576163, 256.6798303961818, 257.3319090630518, 257.9118248409154, 258.26871349423965, 258.5556746618551, 259.1148304673353, NaN, NaN, 112.73099494359683, 110.01179794651509, 108.53793004444258, 107.87087224825515, 107.57119165224246, 107.41565038913846, 107.26075719460617, 107.2514216016249, 107.23692842279641, 107.37033767215877, 108.25663560732075, 110.46963351017385, 113.2614536819786, 115.46268869023869, 118.27482914947673, 121.5298888693326, 123.17803968918172, 124.06825004663547, 123.85198355203279, 117.08031839530845, 114.6981276680912, 115.47231850369892, 117.4560471052526, 121.32130537372156, 125.51714043477122, 131.3892719058768, 136.909389514647, 147.95135683105374, 160.67543762388567, 172.60606802013984, 182.46313219003423, 191.08658734341364, 199.11518636590841, 205.0546095979847, 209.73994716861768, 216.43979001891142, 223.312908299924, 234.42158647001744, 243.39282559525972, 249.35103211898934, 251.90756305568598, 252.31980574363163, 251.96409391469183, 252.79347922293576, 254.58358850052423, 255.88420279399364, 257.97236992939906, NaN, NaN, 109.38974595403758, 107.34054209399969, 106.61116641855894, 106.48135115404105, 106.67546040849952, 106.89027706178668, 107.06638802380294, 107.20523922813028, 107.30150411446276, 107.32416492094185, 107.34975964980768, 107.37534817804848, 107.32581712796839, 107.57373365687917, 108.59960382695475, 109.39594057267547, 111.33857188702969, 113.53341745094298, 115.03032092100749, 117.75699594898506, 120.60577620471211, 121.7080157984344, 117.47636867257019, 116.16995130687931, 116.95394608570457, 120.59588877000014, 123.78562864560152, 127.31606715720888, 133.0805885413976, 138.50388039276822, 150.2416429736878, 162.05129456572277, 172.20730162829565, 181.16614615375082, 191.10914356698333, 199.68535371069254, 204.73882594617362, 208.90499204234507, 217.06913473632784, 223.36844858459045, 233.56214653884754, 241.0071190231874, 245.93303518106424, 248.64406876198296, 251.15034236262264, 253.16862109971174, 254.56267822448999, 256.6284511925265, 258.55236630018317, 260.0386231244627, NaN, NaN, 106.52601479625586, 104.94637756498639, 104.58570923297624, 104.96015680452618, 105.58747318989283, 106.02848219456982, 106.8089612598652, 107.86827562437895, 108.69876072934272, 109.12373583200531, 109.44097838212186, 109.79723870939199, 110.11041817415772, 110.76165302630926, 112.67551849722712, 115.34775066780365, 117.36044474480978, 118.62843768341047, 119.68169272701522, 120.8461555944369, 121.31437051065663, 121.6425212044924, 119.37020844651171, 118.93793441136584, 119.27525211256577, 119.61045035834712, 121.49144864441159, 124.36652185735012, 127.67726710781277, 134.67866458371623, 142.32502223316993, 150.61285591049264, 162.43558090967176, 173.81393205955908, 183.6597961078815, 192.4563768395635, 201.96604784204084, 209.81617202470332, 217.0456376607813, 221.56339192528523, 224.45947680902663, 233.88078615312347, 240.4551588375848, 244.65049211980477, 247.06486285114528, 248.68512705559357, 250.3883917001428, 251.723376858614, 254.1962281725359, 258.6772217618482, 260.82153179921227, 261.9465300951196, NaN, NaN, 103.48226082221446, 102.60948033202733, 102.8696727311279, 103.57404263293611, 104.79673138449888, 105.78581439398016, 106.40471858615888, 106.76392573710409, 106.96981556145757, 107.03019414865297, 107.12899734518021, 107.15482433039388, 107.29001038654535, 108.0561052762158, 109.84002547938735, 111.34490474923089, 113.42975662369348, 114.23895069022534, 114.31531859324616, 114.42416526959225, 115.02159147319884, 116.71098803426092, 119.49114000601521, 121.0374225601355, 121.68946465471727, 121.91855538502764, 120.9591650503785, 120.75605049829441, 121.64282031777148, 124.98230647369626, 132.87747613034284, 139.9506327032809, 144.68576399025858, 147.65383126077353, 150.9640925476882, 162.3750934533773, 175.85678437031314, 186.73702040621563, 196.41612920609026, 204.92140674815494, 213.84452012452314, 220.9652887271316, 224.32663503840664, 226.79864958198888, 230.06126907658586, 234.08572743805072, 241.4315691415812, 245.924662500999, 248.27226350757522, 250.87626549239832, 257.1016561887221, 259.1907467445638, 263.6293351807798, 265.984805329471, 267.3000156477983, 267.15696344324715, NaN, NaN, 105.04410174807158, 103.98471201200752, 103.53780170169438, 103.613172486678, 103.86503803752575, 104.0430989563477, 104.18345935639137, 104.54791742162381, 105.47629283557755, 106.25335809200757, 106.73209658489789, 106.8876544030589, 107.10334942681466, 107.31927692712641, 107.64812208359874, 108.30027227298675, 110.03402536340639, 112.23065838209244, 114.4356311092534, 116.1677476019874, 116.87817353761876, 118.24113799376357, 119.69315812223864, 121.03185234316047, 120.29835371349739, 119.54695768632742, 119.6603874681319, 120.43417257956317, 123.76691134064093, 128.74987999572159, 132.51016906746375, 138.1580277170051, 145.9197469507298, 150.42942523796413, 152.3969539609938, 152.8156837654968, 154.69349925225123, 165.47111115005546, 176.64645996578847, 187.26214509998084, 197.24803762052395, 204.6952134038857, 211.46444501595292, 217.91725193018567, 224.95326893715315, 228.68278358037682, 231.6299911448472, 237.07718588859072, 239.71511424450932, 243.44436253810187, 248.93711353199214, 255.34393817776603, 259.43281053486163, 264.9411811713141, 268.1012455648407, 269.0621247755471, NaN, NaN, 108.01471055552315, 105.13108890845145, 104.14069188021644, 103.99205286802786, 104.17331791490852, 104.8704371792886, 105.9742045838576, 106.89236315007541, 107.74175001319884, 108.69804586100551, 109.65194978075363, 111.31130643644343, 113.78816424303204, 116.38631606196213, 119.091730544138, 122.8638698676164, 125.07122446343034, 126.38135216471666, 125.97458870817162, 124.32270781618465, 122.48161334969413, 120.4418062331894, 119.10699798655641, 119.10403424314282, 119.5522816334558, 120.72969772257812, 121.31928244412245, 122.93583757906255, 125.46158940737125, 127.95885898004529, 131.18920246630765, 143.48134967193266, 157.68937102526266, 168.31159684939215, 178.51773945117304, 186.3391295978755, 192.82243893814217, 197.9800822848354, 204.5669605741916, 210.67197481539154, 216.5919705403049, 225.2589028208721, 230.9499366255863, 234.55947689718099, 238.47638307103423, 243.08338275309768, 246.35861456092613, 248.81597084666646, 250.89824687938076, 251.6491352311528, 253.73310158423905, 259.286338787668, 266.72857817414763, 269.2939391109898, 271.30960271231777, 270.674059451828, NaN, NaN, 107.04484646031796, 103.4091045094952, 101.75861689781394, 101.46752103426178, 101.72324963980329, 102.5681658298551, 103.1524400879294, 103.58605064542841, 104.39043230290189, 105.15644181850536, 106.49021320981683, 107.96922884730522, 110.55493005459354, 113.3486933932963, 116.22767686657244, 118.9877904309523, 120.93392517048375, 121.94949196797764, 123.50494898543727, 126.01647740136791, 128.21553137068605, 129.66960443669808, 131.5741776164995, 132.60939289930485, 133.07936143385237, 133.95526806394406, 133.65770349245793, 132.51239240865738, 129.29819639936068, 126.35749900853395, 125.49376608505395, 126.52486896119129, 129.47810172431915, 139.40522751583873, 155.8213919963297, 167.19840117868284, 175.46860567328966, 183.14904795327382, 191.4591115687717, 200.9855104291662, 209.274320667388, 217.67594825594782, 225.49838460696247, 234.66098901130374, 240.0452432816922, 244.0740825719766, 247.995708020247, 251.5466286575425, 252.46824071415193, 253.7290374258416, 255.1341064139688, 255.03723845704036, 256.7497862358256, 260.2424461464036, 262.51072715390893, 264.10549713605485, 265.45592103405346, 267.37689254214376, 268.2543437941985, 267.4077843540301, NaN, NaN, 106.33810281288467, 102.29738422138828, 100.52901697669549, 99.94069457978762, 99.86224012891813, 100.07755967621196, 100.29218166971529, 100.57976644830329, 100.86556689352986, 101.53076173535108, 102.554244044, 104.32229384249113, 106.31326046612588, 107.92774264391946, 109.77570083526709, 112.27457652448753, 117.21061575700466, 124.11205973388627, 129.31992844793615, 132.98023699558027, 135.5849090773028, 139.4166373673337, 144.56932484604485, 146.03540063254425, 141.20329200658884, 138.01526103113008, 136.586709520346, 136.31978712341038, 133.39814903744642, 129.00897032542096, 127.8457061594847, 129.62008562325335, 141.95490477888657, 159.26493833575168, 171.37430235353696, 177.84971902560096, 182.41586965898347, 187.43907634226602, 191.5585229580141, 195.0985779627471, 197.53581970393805, 198.92432625600227, 201.7418365228805, 207.21478781465697, 211.88965677659405, 216.17628749580626, 221.50078722497406, 225.573368639939, 230.771862407705, 237.5476549889654, 241.97474633471333, 245.93664653533062, 248.78690908448573, 250.1613154946225, 256.2583531643131, 260.12111155341313, 262.78362564269776, 264.4551952177579, 266.2121414534832, 266.7802967397919, 267.5740631374774, 267.85518523679315, NaN, NaN, 115.94390721790823, 107.4986240444334, 103.16609407101434, 101.39979775285282, 100.58616658414405, 100.36184993897731, 100.42870400137188, 100.64133179423872, 100.9268031962589, 101.2148091663696, 101.58177156268344, 102.53232545965331, 103.4803690952363, 104.65224016037851, 105.90102382675705, 107.44365201027792, 108.84013463576329, 112.5173466054006, 118.01600282432236, 122.04224158250445, 124.23752461816655, 126.1367687581258, 131.42568494401587, 137.17194513188232, 142.03502562150848, 145.5722703137022, 150.75668211958254, 154.41769773180633, 151.18950518175816, 144.21311861889532, 141.5934815802412, 140.44297615497706, 141.63570635714163, 141.06421278403212, 142.8637708593378, 157.6965808863808, 169.1931775841621, 175.6658160596743, 179.17971745019247, 181.67264010295906, 187.65633417860775, 192.5928270020808, 195.46132148520826, 197.76388867040745, 202.32569040929243, 209.1421032693893, 215.27719891902072, 221.9854296623253, 231.95363950012398, 240.74539501927165, 246.13295281059132, 250.0108689353359, 251.26810558176695, 253.0765791782972, 256.7807034574487, 257.7444777105248, 260.78590323603356, 263.70631517077646, 265.508449999515, 266.7868518246224, 268.1866545429503, 268.82150749990996, NaN, NaN, 115.99140286790941, 107.02963150359027, 102.76350272045913, 100.55724335707374, 99.59721063639464, 99.15098207567861, 99.07130591102398, 98.99132722436876, 99.12303395267266, 99.10968206571246, 99.17385895270132, 99.45715909609076, 100.18574921148273, 101.21132487729147, 102.89985718587356, 103.91442387961793, 104.34226156333561, 105.22267030038905, 106.69553646969558, 107.78963066040926, 110.4344118217136, 113.4389332181506, 115.92144309313547, 118.7012742689284, 122.66044558606994, 128.4650674462463, 132.1616811206254, 134.60897576113481, 139.031383684813, 144.1147471829426, 149.48521716653119, 155.08952129355418, 159.7101189970469, 155.17317422474238, 148.45861350995693, 145.83828492473148, 144.73977285207064, 144.82065071582943, 146.64124983265455, 149.61567200962088, 159.99148423192554, 167.93330122770456, 172.8966751643383, 176.42601117172674, 180.29781344346702, 184.9797981297708, 192.09549997733876, 199.03727387100983, 206.81824470193848, 211.9023678920603, 216.7143579446531, 225.09720205100072, 235.88180443703078, 244.23986218043927, 248.696473667374, 250.96308841005305, 253.0665211314637, 254.4861864255088, 255.3169186043999, 255.9636418243775, 257.09600611968307, 257.7417652684416, 260.61503990831324, 263.96120146997424, 265.9881079886476, 266.11189651603644, NaN, NaN, 96.26674341755611, 93.721909287246, 93.15895472525185, 93.03568742537087, 93.3465744697275, 94.21423147245861, 95.29679384684611, 95.93796315847072, 96.57856823597389, 97.77564400334013, 99.75169351701062, 100.84045485329861, 102.8199030224902, 103.89798121213424, 107.53403302491728, 115.22575870589608, 125.367515162293, 133.00441649101657, 142.72588635322145, 152.13813067250575, 161.8982095508012, 160.68032432682796, 156.84874599894619, 164.3975099193192, 172.95242792233324, 179.58987978958257, 193.1961682063387, 208.27914578702718, 218.64024860117107, 224.9939527254715, 238.25183136726156, 245.70651745338407, 252.22792672924922, 254.27544077945737, 255.21697846737166, 258.198420290884, 263.78746566108686, 266.90845621578967, 268.20629964585777, NaN, NaN, 79.41072607237722, 75.23688850330771, 76.68459129186138, 79.89368733760568, 86.62274629958108, 90.36453715476583, 92.88651159401014, 94.96965927175673, 96.39047436334785, 97.92030787098412, 99.22722624668008, 100.75607964833995, 103.16468767994944, 106.13586449558925, 113.38596445913493, 120.86134747455716, 126.4917983651122, 132.69828221716554, 143.2345754154161, 152.7449209831532, 159.8671532355274, 167.6737830211109, 174.49084953349856, 169.52081863845564, 160.01758409192783, 159.00369730516312, 166.23760613433268, 174.77659136490928, 184.82602502255017, 193.16061432716015, 204.8755216745277, 219.76262377925946, 233.549563725452, 244.1844072637583, 250.79958130117785, 252.89485637559181, 254.81070389580668, 258.3416104301552, 263.0546509713212, 266.2069232256417, NaN, NaN, 73.31036829573497, 70.88451752376639, 70.24772149476456, 70.16225971964548, 72.1480855022238, 74.12182815974205, 77.20763929053138, 81.28519622160753, 84.69273670545144, 88.10448697273844, 90.07248510238323, 91.15681850655032, 92.46645326206844, 94.43639195239871, 98.27103650157923, 110.26242421082964, 120.50124626574377, 124.37494737432117, 124.93770430869547, 124.63219079255653, 129.85986524229412, 136.51063606707004, 140.34489991946728, 139.31565762379145, 137.41235792914554, 142.27665394608974, 143.61567430830743, 153.96805014146776, 167.5299226301377, 177.9851403409995, 183.1610936786669, 177.20862062504784, 178.9606431862116, 184.5632453829379, 189.05031032916438, 195.9878519763737, 213.13678922823297, 227.5574116581601, 238.07139479889713, 245.21430295484214, 249.95115021307936, 252.16456344315154, 252.91983860492388, 259.9307432500334, 264.69040720465244, NaN, NaN, 69.50913311603743, 68.76792085024275, 69.05272085057153, 69.33587547300438, 69.90749751397692, 70.62702466948532, 70.61106771276758, 70.59638782968392, 70.73498210190235, 72.81111848222471, 74.72259310483476, 74.14061131068769, 73.72387680730941, 77.55947194361933, 80.05163100407238, 82.25827189606446, 86.08195686835023, 94.44221967946734, 109.39454647165267, 116.89129313617163, 119.53789423276577, 119.89344084529313, 119.86279331007864, 119.28820392167346, 118.89974973162013, 117.9801142350594, 118.14764636130224, 120.18232681113089, 120.40177629790301, 120.93769123868549, 124.99917364974536, 134.75656481182483, 141.15209686457752, 143.3319645598028, 145.00865940848024, 144.48402147486905, 140.15220932472667, 152.74207050507283, 175.1098133893624, 184.64340498153456, 188.88251905342352, 193.62492284666345, 204.93827808392788, 217.19418062107096, 225.09771471703638, 233.3304600579144, 241.97178182796813, 247.4872557532294, 254.27474648296678, 258.0717766510572, 262.84232059574975, 264.4755623697718, 265.41479230246193, 265.8171322034393, NaN, NaN, 71.22259033602337, 70.19152978778942, 70.63045492035465, 70.92423678065718, 71.50838533452121, 72.53697836998205, 73.7151919001167, 74.8879421835776, 75.7645929629475, 76.0474673667132, 75.75011436557566, 76.33753235908121, 77.8162356516109, 82.94823714960377, 88.21838100188896, 89.96988265909077, 89.81732208080523, 105.37784264999041, 116.81136970205269, 121.92953274097684, 124.36268493028996, 125.10952919781616, 124.24488858131065, 121.1766527742921, 120.28335668017277, 126.33925675413361, 135.71221251690974, 141.9045938782831, 145.87244855518233, 149.1934595777436, 152.4159562538494, 153.9021571671246, 151.2167481655378, 148.0146514171195, 145.9390882681914, 146.279636971176, 149.57665744665684, 162.19297087643665, 174.82143033527802, 186.31726079484497, 193.52711174486188, 202.2569330305705, 208.75162734988652, 216.9404398819535, 234.11046234276267, 245.48090141049573, 249.53659183082624, 255.44292950196265, 261.1199763096162, 263.8353814555559, 266.4594156297465, 267.07182678920736, NaN, NaN, 71.3778557659611, 70.3419710446792, 70.18883486810692, 70.62603820413584, 70.90915835917126, 70.01463545694814, 69.56665185591555, 69.70357483131687, 69.70021180555212, 70.87755549994145, 72.35009490722092, 72.48053631455505, 72.3209388689341, 72.46094106307672, 73.92581551405252, 75.9803240551655, 77.44717580346794, 80.08395346750359, 91.98193917288562, 106.49954000990702, 119.10413287831172, 124.10385781803548, 123.15731997915414, 118.24948823354072, 114.19524006211081, 111.83334499777425, 120.92639767839941, 127.67351683419358, 131.86392386616293, 135.76101095684467, 137.27518067774014, 138.211980125135, 140.72346714395673, 142.60933484942598, 145.59387459865948, 151.49761214253041, 143.84113161657768, 136.1387500308597, 134.08277752998364, 135.84636128989828, 137.8547704205387, 140.25211364874485, 142.83459915602722, 144.48412573614007, 147.07344033357984, 150.5818733693112, 162.07931381100383, 184.67835296393295, 198.62174361907762, 208.89600397394005, 216.1686968370473, 220.09707308686797, 230.97557713080718, 245.1101802446746, 253.35096226254677, 259.45841425825887, 262.25604568573584, 263.7051352849615, 263.75618109548765, 265.8502057596973, 266.3428365865725, NaN, NaN, 63.22241629620226, 61.781696032533446, 61.961711599451625, 63.50831648404209, 65.27324291907343, 66.85284779145655, 68.27713022107305, 68.88752895320589, 69.13157229653882, 69.30250225315447, 69.54499976148992, 69.71485553946418, 70.18187903233819, 70.9827666531592, 71.59815006619698, 71.9206804304918, 71.80079504375468, 71.29112171911726, 71.0216630518774, 71.00503501486563, 71.33507420542207, 71.62321461228798, 81.46424385591187, 99.06584573029329, 103.88851152686578, 104.31014351714755, 113.25618230583397, 125.13391523089618, 131.28280985116822, 132.1507225502619, 132.30271632699504, 132.1579447293208, 127.9228742662675, 120.45929766859457, 112.38393953715983, 115.61778662792898, 125.47890869476869, 130.9195472489254, 134.4490940704976, 136.3396227836384, 138.45120682247975, 139.58531510135387, 141.8000046377779, 144.21157782901608, 147.3660865266538, 150.75818252370118, 141.84152709991486, 138.69346941334513, 138.86348038459764, 140.5237041700842, 141.9828777707345, 142.6987842671292, 144.35549568609463, 148.063054860085, 153.0466661608824, 159.7539248854109, 179.512342894096, 195.1368570489717, 204.93943030079512, 212.67293867176355, 224.31637642251363, 230.91656030822577, 238.3449504043159, 248.75487936604787, 255.87601702367328, 261.80392898607494, 263.807883468539, 265.1444304855034, 264.89005632795687, 266.5711178516331, 268.1818466138147, NaN, NaN, 47.47985761609835, 46.743948042180236, 48.03749913155742, 49.287152964837375, 49.71681180461418, 49.81575830731694, 50.099900445374566, 50.49513011919065, 51.26001982389667, 52.83927050980055, 55.006893995412874, 57.174433212284356, 59.15465521238644, 60.578622520093425, 62.447390277661334, 64.31516992664977, 65.62636913520842, 67.6811889385653, 69.29924176040777, 69.8020129195561, 69.79767644237319, 69.3460902720782, 68.89222362094168, 68.22177849298097, 68.65438445463805, 69.30203952186406, 69.5145825187423, 69.06209131779943, 69.49439803597642, 74.34610065345248, 78.97119318704213, 102.74692274573835, 117.70507846786192, 124.51884942028582, 129.36016693157654, 123.8591816865357, 112.83879706360845, 105.57552001370814, 91.49609977295606, 91.70582141133086, 108.65216934470044, 118.90588120061233, 123.74441479565058, 127.51593529426253, 132.74031258810268, 137.52798916240172, 138.506105795282, 138.83332532645085, 144.3662235444092, 150.88360949649422, 158.28960359521093, 159.5136973909879, 158.87711674446808, 160.00433859401215, 157.13453310857972, 152.76317330266855, 159.26633642177487, 165.5523611738907, 169.04407515741792, 167.67414497603656, 176.03669820411082, 194.41828817954902, 202.42960349907494, 208.2921032774801, 216.99574433417408, 225.09732098048627, 235.52643822055074, 242.0631643333239, 249.58210457083328, 257.4764840556736, 264.0954383922505, 265.6889512375087, 265.6202022593208, 267.1591969063148, 268.206508118807, 269.1507661445873, 268.79442932781365, NaN, NaN, 39.49337781926027, 37.355479022025825, 38.28491108206891, 40.78532124762286, 43.39611943286698, 45.306665539933846, 48.39299599779507, 50.9340462131992, 52.767145821254324, 54.08458950317921, 55.85089147840021, 58.5716580610669, 61.027644091038326, 62.856014622742535, 64.61123985093394, 66.14734763210524, 67.71969777565839, 68.70091579837106, 68.63723551531143, 68.55339439072898, 67.70965707649925, 65.39280259785913, 62.84771391835819, 60.743528435019, 59.52163004423086, 62.27174022973787, 66.34530040400034, 71.95769747396615, 76.57883469068742, 78.88782348242611, 76.91178909878442, 71.83545977586392, 69.06904830734663, 69.1664643207305, 71.13470621828316, 80.4772464731144, 90.14636790519302, 97.17543115222774, 102.22487795948092, 105.40462926811202, 107.6333353893193, 110.04316637410257, 112.79580037405172, 116.54375878594846, 120.41042343674873, 124.52640148042137, 125.95203184783774, 128.59610078359853, 131.02714674204114, 127.75581999717247, 130.5145277756194, 142.13672984635022, 146.54134469168406, 150.4077128154971, 158.345769691057, 165.34607313284727, 167.58962196554106, 165.717961966027, 163.5430989414307, 162.23708161746256, 162.39541947609644, 164.74625896677247, 169.05735383360658, 178.26248216074538, 185.9201370887537, 189.04992638746077, 201.03393704583257, 204.195134396686, 211.7799640838609, 221.07014900735473, 231.49282977310088, 244.39940872184377, 251.09184104712511, 256.2817225319457, 262.94713870103453, 265.2513479377608, 266.01752788751634, 266.511964589571, 268.0500015484743, 269.26393700600255, 269.7235510539246, NaN, NaN, 52.797179204792315, 51.94543487499853, 51.75890075033062, 51.78859362938588, 52.19288530641733, 52.85118213594936, 54.09931607727348, 56.15470923274389, 57.765635766675366, 59.52496183076014, 61.13465273813506, 64.2267774320138, 66.83107390502065, 67.85164136721285, 68.33295053569907, 67.15612418097639, 64.68851522966546, 62.473900838487076, 60.918738016971766, 60.06090426659679, 59.13194204356493, 58.02239022360978, 57.64996325463424, 57.055770193591165, 56.902238045326754, 57.03784840352464, 57.10225073645752, 57.389975949493554, 58.48352350031773, 63.46889616183862, 67.42725236670186, 69.25377924393892, 72.55333727928605, 74.38187616602725, 74.37668764137275, 72.60451039979623, 72.97253503073932, 70.98137015210325, 72.95366500373181, 78.0110139858676, 92.818180418575, 108.53161555677445, 114.98616558973318, 117.92069631032807, 120.1033624389603, 121.8591539303053, 124.8209033699643, 127.61396926702906, 129.8127307127626, 131.72007107535018, 134.67723351554235, 136.7444351062635, 136.46036935843966, 140.4619000539173, 147.09656482023058, 151.57313941921518, 155.8689221998117, 157.34212124122425, 156.21320153498607, 157.48224336349196, 162.09795719673912, 167.57145285567142, 174.83993865322608, 182.404159236105, 187.66778534198536, 193.4997209828918, 197.99715483985133, 201.7895290380969, 207.36646539754759, 222.91545549406052, 238.9246272640737, 253.6415518466959, 262.87088475974616, 266.0277874640898, 267.68965940232107, 267.32872422124296, 268.86789063935765, 269.721540565345, 270.7204061304236, 271.2145485245848, NaN, NaN, 45.86583529627752, 44.57293900248208, 44.4974185901306, 45.52756408072908, 47.76732804764206, 50.04727580486576, 52.36698661770806, 54.365020483506, 55.75351391262989, 56.737231759304095, 59.749639505440214, 62.875787152153706, 64.26768574120693, 64.55196367529905, 65.09727186562145, 66.34024719741132, 68.15031999497383, 68.36568755349721, 67.80066289206879, 66.83423702667858, 63.89108892165605, 59.76936192501354, 58.436860638388694, 60.34508355147762, 62.69130332950848, 65.03709110100681, 68.26096299956822, 70.3052277931456, 74.6994883561518, 80.41454130908933, 88.18586509657592, 96.83855414367207, 109.16529744065173, 117.3714278005323, 122.79148012692914, 115.4654020689123, 109.30516046617402, 107.84081284311182, 93.16597213577228, 83.01674917714313, 81.2402141519806, 81.77916932199003, 84.18960510952381, 88.03380228865022, 95.07987692685455, 103.66100194399323, 114.98525318263641, 120.70065384263245, 122.8039435423783, 127.9771355831142, 129.8444218553928, 129.8415534167836, 130.2079468068899, 130.99605956878062, 135.33555631716806, 142.32789835683656, 147.77966774911528, 150.39548835951265, 150.1270241979584, 154.1504363235627, 158.16183772772553, 163.89697729704517, 169.6176380691031, 175.55007318868368, 183.90403838615885, 194.49573681905014, 199.1852195709011, 202.11523657754188, 209.10408117092712, 228.68873201017828, 239.27890563083085, 249.11884821420176, 256.159956554932, 259.3273816847632, 264.143375723516, 266.9348824477411, 268.486534130325, 271.0579812311835, 272.1982742437278, 271.914403556708, 272.07780391292863, NaN, NaN, 52.03366033644726, 51.29174155346312, 51.211310104731375, 51.424646300847044, 52.19059077988667, 53.065211221546335, 54.1246431752365, 55.44657148092778, 57.20872233920153, 60.269516381220946, 62.6574889907781, 64.1571891055957, 65.10333000448544, 65.71575953024562, 66.07261885435724, 66.65049438619624, 67.5609022486621, 68.39902592149222, 69.09575826539863, 69.05146860877792, 66.41047237640137, 63.281740102525916, 62.54176182937249, 65.65711760866257, 69.14168196303586, 68.58799541676787, 68.02506179466437, 68.74782157299154, 70.39124492667767, 71.66779854594536, 72.39403743541172, 72.02284145547893, 71.27800762829307, 71.0867936069025, 71.26972572731412, 71.81106958032282, 74.18918904355137, 89.77838753481369, 112.69627367045914, 126.63913200101862, 131.70177497319446, 129.49401949484155, 123.54014607151457, 123.53435680640241, 123.74834243649155, 122.63931048561402, 124.3950697211501, 125.49029500039708, 125.39190670610476, 124.95569354383836, 121.35392269495465, 120.81191093296931, 118.95977269016016, 118.08162994763578, 118.52562278539023, 121.7291867842371, 128.56973873845698, 140.95017690735102, 144.05004297954153, 148.73797169670428, 152.01786434423107, 153.06423753071428, 154.08552412251646, 157.35766965276167, 162.46561954413505, 174.66102694242642, 190.3493251697481, 197.9624829681489, 203.3692422476589, 207.13210478017598, 214.46516751952018, 223.42429932111912, 232.49314813391996, 240.51794325934728, 250.5390234184389, 253.59490844265372, 256.7762617760499, 261.0423040972107, 264.79800431681883, 268.4380300178694, 269.99813192884534, 271.1229601631956, 271.031613233494, 271.54008070641424, NaN, NaN, 55.019633884971796, 52.0677886057115, 51.65814435399553, 51.835408860259605, 52.15705488598648, 52.48095116722946, 52.8782491004519, 53.64808714781484, 55.04008455875388, 56.68780534731998, 58.262806127668696, 60.65316599112469, 62.076376627980764, 62.762475483652814, 63.970751004313506, 65.88563706739296, 67.90349348771238, 68.70324608755163, 68.58811670431051, 67.45435665846053, 66.23389700605382, 68.24855370813512, 69.60085770734962, 69.15000926538598, 69.35919626847243, 70.0820392298036, 71.43148220299452, 71.38423939249813, 71.29996312956433, 71.10530109411967, 71.16900512280552, 71.33823666136973, 71.25624535883217, 71.7982883213202, 72.62891398019752, 73.94808992206379, 76.807684347868, 81.06942547399309, 79.75090564963043, 79.66767449444458, 87.46610286715821, 91.85522322180364, 96.24928708958619, 95.14440225162787, 97.21901830641903, 104.35783716542994, 111.1702870819098, 119.31442946481567, 124.82136566156547, 127.83091401989064, 130.81258656804337, 129.7253567773314, 127.33803735089273, 133.9875029449732, 146.5041205226754, 159.40436637059608, 166.15852404394207, 170.5800029073861, 173.44053483911307, 181.26762439256214, 188.03520275444467, 194.8891745913274, 200.17297041710486, 202.7761956506202, 206.20355728252997, 218.06261652639876, 230.22053529065582, 243.34925951665232, 248.93108003605903, 251.8941371564927, 254.42521032038871, 256.68669000703665, 259.5321698736966, 265.19679632983474, 267.3037091391497, 267.2015870664528, 267.66634414272085, 267.6182563156523, 267.31369909021936, 267.37902226322603, NaN, NaN, 40.653741168719826, 39.50926772377099, 39.61726220446887, 41.35006384443345, 43.73963253686589, 45.53921028109964, 48.29920450123132, 50.27951372569784, 51.92988493618356, 54.764149083249784, 57.37610860340874, 58.655972343864974, 59.19964651167296, 59.781193832432855, 60.913855547939924, 62.52337463217271, 65.01746952353807, 66.3654703706687, 67.20051786336211, 67.22961491639606, 67.52230767580491, 68.39876923590533, 68.86893198467594, 68.60330960032215, 68.78919482260993, 67.42446814644832, 65.06803934023927, 60.54914875588593, 58.33856929075026, 57.85232592425023, 58.80028875385867, 60.517679765443106, 63.66868652724456, 67.81503365227759, 72.28985166414513, 71.26011543485468, 71.18900581398658, 71.32820402638241, 71.53539600730632, 72.41007865839134, 75.45683921810664, 77.2099657759981, 77.53127354832597, 77.8552162698579, 78.40195826680436, 78.2875660450247, 78.3909310546471, 79.04049031391794, 81.1179164674864, 81.54229028571744, 82.2993784448756, 91.86199215932633, 99.33384743674382, 100.53031401930171, 104.47715481270887, 107.11309703871932, 108.87319890230893, 121.40203172053155, 127.24123757478021, 130.35968273116194, 132.94736675189233, 138.57096461025975, 146.99056715270063, 154.71975687335032, 162.7599813911788, 174.16473594395845, 182.94100749214272, 189.35763381408043, 193.37719393562065, 195.41770658807255, 196.5593969642798, 202.88685875162773, 217.38289065361155, 230.30781341707646, 242.6349338135312, 246.7511300647253, 250.2137843809886, 257.6673464332885, 265.5471571243761, 266.46863079144464, 266.68002315759645, 268.15573027433874, 270.3843353353303, 270.88613518148657, 270.3948292450421, 270.61272329831564, 270.88572917971555, 270.9609686949672, 271.04732181917035, NaN, NaN, 40.94575851111338, 40.17092538263076, 40.68391553936063, 42.26709788624709, 43.50898929557927, 43.93988629009959, 44.2603807144657, 44.987434476357095, 46.638713017804214, 48.72891342904249, 50.41440745683658, 53.06020471320732, 55.04136766212778, 56.76316974177193, 58.59993074269173, 61.39037319606757, 62.590148531278544, 63.09216913654814, 63.816436200149674, 65.9140048830283, 68.15419883410789, 69.24842163728975, 69.50917091901864, 67.8949866671694, 64.03682866852134, 60.58886190700549, 60.39673281344096, 61.89961977919979, 64.76288686422332, 68.43584659549205, 70.9358732704924, 73.77295239160676, 75.12017619541862, 75.58653744857905, 76.2080740806304, 75.83594859567563, 76.79658046963216, 78.37849810417922, 79.21733888625504, 79.6515227901597, 79.49651189707107, 77.50749809092198, 76.91291427737201, 77.05254928253524, 77.41164994070576, 79.68650900049303, 84.31285895064202, 87.3848808499119, 90.47179330188116, 94.65782928043714, 98.18811496311977, 101.71685334939782, 104.57119520413747, 108.7526806834947, 113.62153951707327, 117.38360037548732, 120.40516400472525, 126.64355665253255, 134.87959059455193, 140.12823498079266, 147.0417946540378, 157.05838220161687, 160.3753268552732, 161.1557888778547, 166.64846998882055, 175.38983886828163, 181.580435113927, 187.940097230779, 191.93387763442357, 190.19612426281827, 184.32852987371658, 183.43255412661006, 186.84617999915162, 192.63846478065065, 201.2591380572215, 216.1672415265614, 228.49023158463783, 239.3707938413829, 244.69656709844597, 248.0564757710401, 254.5728352214402, 263.11858130230263, 266.08369600232265, 267.2717562988627, 268.35829192513575, 269.1779359557189, 268.92007948448895, 269.504137769212, NaN, NaN, 45.27039868919937, 44.38511171675503, 46.00407803622888, 47.83577090432525, 48.63530517205669, 49.877637881800815, 52.30584946848507, 60.575611784504304, 65.87145520211217, 67.03278617581755, 67.23885453534008, 67.3716538506863, 67.65100506710759, 68.0055957791085, 68.8087735754142, 69.31553496157153, 68.86429987807765, 68.1185245912533, 68.10762180063227, 66.85536108551673, 64.17228385720921, 63.73371637391806, 66.22749197381393, 68.0524024512341, 69.44449982914786, 70.99634556369472, 73.35312012352522, 76.81717317137667, 78.8654047295933, 80.11484735133682, 78.86541529829265, 76.95047583254166, 76.79043993362966, 77.07205359301628, 78.31292704755806, 82.3558463546177, 87.12842466160349, 90.57336083900648, 92.54062945152052, 94.06582610853994, 95.11445925124154, 97.97673667703074, 101.82752302254413, 104.33487021470408, 112.04959277029475, 119.21969806149181, 118.36386198929497, 113.8495101603464, 116.1023309277206, 122.8430100878211, 125.71153331012808, 130.91866880366226, 140.02029555254654, 153.14401441292725, 167.0067763690144, 178.0108595000351, 185.20951552970934, 183.2273251332341, 185.66648199859893, 194.90248471552047, 207.98002944278417, 227.8939331007215, 239.26799150224986, 245.84876130722006, 251.5549005252071, 257.6178064412035, 260.5667180272923, 264.6745991944294, 268.29384833353225, 268.1256467542332, 265.5447838899276, NaN, NaN, 69.30725543409457, 66.86976459355759, 66.85592014820587, 67.27354553489351, 66.83788227010172, 66.58642009296493, 68.2357134836978, 70.40247412396218, 73.19874186433421, 77.09499842539215, 80.21883830739546, 81.63655826779892, 79.96902367641377, 82.27635417287189, 86.53082429820009, 90.22664818792609, 92.55828222793208, 95.47227630647875, 98.64147009069194, 100.04865385555337, 105.02337019783941, 112.50084950464176, 125.73034867820209, 132.10186391731835, 135.6066974391272, 131.06554253569573, 123.6698372947803, 130.0940595637875, 133.60588397809926, 138.92886467041347, 144.91590729075733, 155.83098783338443, 163.57485607557848, 171.59239418667585, 191.1569817102581, 215.39609315141033, 231.49888836068715, 242.38314848274757, 250.8887286893237, 255.30236453655905, 263.8039312328304, 268.9731199023399, 268.8267803850251, 266.33008049624726, NaN, NaN, 78.664791724928, 79.99123641924821, 81.16923132363668, 81.90164639078759, 83.9503007721373, 86.58207640278427, 88.4730295914032, 90.66088488897272, 92.84430143817518, 95.1755695125783, 98.09230813416477, 99.82213844678063, 100.08041238963611, 106.66816468569462, 121.9429647870585, 126.46789142013269, 128.64021605365198, 135.72021558514663, 128.9558102546248, 134.76965375442182, 146.64207362978368, 170.42337390682786, 204.21335186346434, 230.42563638134257, 241.53183650437066, 247.25375076203335, 249.8389071537575, 259.887486718566, 267.0052566548556, 269.1829446069718, 266.8418303480477, NaN, NaN, 91.27057976070336, 91.78305723126407, 93.5709618430051, 94.82894094095549, 95.56841885158966, 96.3035155637225, 99.86636576357928, 103.94961845997443, 106.7467207597304, 108.0075331904507, 117.76932207060746, 124.2103332814354, 134.76664494877897, 136.12010972918262, 127.17740191185923, 139.10368763928474, 153.329716037982, 167.62314678846175, 199.03511678028295, 225.54771489997125, 238.69359476892132, 245.41880076165353, 251.0945583694106, 262.0526710356059, 266.9907490496769, 267.7460581857068, 266.8992957089131, 265.52498020914595, NaN, NaN, 97.78272292955948, 95.19232265622013, 94.912070299744, 95.1361535552567, 96.90261206422055, 102.53548833761927, 104.56206634081363, 108.13274456821796, 112.98439032051522, 121.48116976359319, 124.83562120315395, 135.11091144514148, 141.34079576354256, 129.34129755867153, 145.13310370943145, 162.2023995259911, 192.38638569153736, 222.77387138364375, 236.69010206870504, 247.1406303312559, 254.9666815505868, 259.30606441529073, 266.56761448354723, 267.67393286961175, 266.5215457093505, NaN, NaN, 97.30071795932469, 95.44680884689731, 95.42407370350101, 95.7578474092301, 96.46236015735498, 97.16571058044369, 99.71047260258727, 104.45345001448486, 108.46396350379202, 117.62347268269531, 122.03792185620037, 126.44225542352378, 138.25103855507373, 130.6350751809528, 148.02937692389037, 178.79556046936037, 221.94216256158165, 239.94013374928764, 249.7922594171982, 254.34813622975776, 261.7733436253824, 266.48900801458666, 267.7063161020396, NaN, NaN, 98.37267236760894, 97.17821849614201, 97.15809012949907, 97.71135384210639, 98.26643395320626, 100.29592186587624, 104.09314816218344, 109.36697208219957, 119.93871660781676, 125.25150529582768, 135.54359218305572, 140.80885706516585, 140.84127350309547, 133.52871623252784, 134.79338417066745, 160.8227662435275, 195.56817186135996, 222.5600494262917, 233.30507999748767, 243.00011411790567, 249.21160111199006, 252.2492853426189, 263.16145959744193, 267.954596084857, 268.9207148842889, NaN, NaN, 101.21602110770952, 99.1399035522867, 99.11687228551038, 99.08127796235046, 99.04624944400017, 99.78072524547197, 103.35778751712327, 110.27671225027476, 120.80521455736252, 124.65850860550022, 138.630272084451, 136.1698439083777, 148.07989212717558, 173.68788655605996, 205.97856696264444, 230.2262743126351, 242.8892570666666, 247.77488330606585, 250.0630159510601, 256.9586166171002, 264.1929781186795, 267.6018484522421, NaN, NaN, 102.16700430959658, 100.09063416209631, 99.80769082289207, 99.76798644328976, 100.24764904146875, 102.52995706815912, 105.58000058478929, 110.69797468244715, 121.51669324266022, 128.99109079559514, 138.85348673619825, 131.75556017696047, 153.70323156388665, 180.93232045286675, 213.48892170266672, 233.37283536764443, 242.5424012481131, 245.35875648367335, 246.86487905931656, 252.76225699887232, 258.989949316709, 263.94183264888613, 267.51842917224207, 266.9456210867613, NaN, NaN, 104.60663957420715, 101.24657208777465, 100.70801825702918, 100.67350536145813, 100.89583790971915, 101.63450880586535, 102.88805206057944, 104.1406386385603, 107.97069705644721, 120.32371155626973, 127.28497051862847, 137.12696051158167, 130.02689084542538, 144.74951155471504, 165.92702763804456, 190.63394110590124, 219.5119368342377, 229.8983763534433, 237.06103950866984, 245.22708254706612, 253.26482888974712, 259.9669006949375, 264.79318649530865, 268.36847686610673, 268.51972556041505, NaN, NaN, 103.95327036721713, 101.73253176723527, 101.48612942635881, 101.45221826865703, 102.29865905915337, 104.69806041731368, 108.434855796611, 119.89618634293699, 125.84560311331946, 133.1721598869376, 124.24626538803373, 137.9748958556036, 153.43239876124895, 180.144512338214, 203.98577041610363, 223.56987906926568, 229.3654443245525, 234.55856042056178, 242.336249806362, 255.16255098498797, 260.99609770312435, 264.41835518250633, 267.28713753998744, 268.98001191133187, NaN, NaN, 103.12196668350174, 102.58938691069505, 102.56519333905301, 103.04829318825568, 105.08242197165644, 108.41013615957209, 114.55030572838548, 123.55912420045647, 130.7983713315454, 125.19968259678062, 120.3928662361093, 130.17462383920787, 146.92274183855795, 174.41217474384644, 206.07339257078198, 224.01908881892967, 231.91451388395484, 244.3531713357145, 255.40781008920632, 262.2022367022328, 266.2733883571222, 269.8102251550056, 268.319933878574, NaN, NaN, 104.98121975996634, 104.37233511842402, 104.64547520919002, 106.08417163369846, 108.11161558849574, 114.85175871841034, 122.75522842333685, 130.7262282871557, 122.60016523101213, 129.130752422712, 147.10372972808548, 178.49977313676257, 211.1400675028376, 234.072977916496, 258.61785381849825, 266.92611793821885, 269.2522102054533, 270.38528415062046, 270.64295184021944, NaN, NaN, 107.85907101938369, 106.38401160848271, 106.18134141805719, 106.88752620041626, 109.98889763537895, 121.56909982960339, 120.92183950409105, 123.93108833933448, 131.99323675099924, 142.85474363588233, 147.78906713525274, 149.24111984063165, 165.3201002609942, 182.8793273457596, 206.30232712458618, 220.4060141804039, 234.6302353890339, 256.05226866050594, 266.18675327492, 267.7238576946492, 269.05954238473316, 268.6279388172807, NaN, NaN, 104.84575924477367, 103.72648363658239, 103.25844287210536, 103.44035969674954, 111.8318639813566, 116.49893046266932, 120.5320726897014, 134.43923810353635, 148.5671303925112, 159.16844585772628, 181.58545314163675, 209.15744626523198, 230.8274999269784, 256.3958761078541, 266.4762877011082, 267.5147885763478, NaN, NaN, 101.68592219432487, 100.12435809688463, 100.09932823846636, 99.84315364420914, 98.49613992463826, 92.97824573376344, 102.22843774800762, 112.44978001313524, 122.38981737644897, 135.61135030482066, 153.5340266269902, 170.3290013784361, 189.91627143211255, 211.47291189157855, 238.43898897645948, 260.63764532796523, 266.18359762354294, NaN, NaN, 94.44685159886234, 92.66567280770843, 92.42241360246948, 91.73570658969672, 93.03881238467551, 112.25350677763409, 108.77150371054832, 118.03494913646088, 127.71624277940045, 133.42125938784662, 148.02056264726522, 164.17084173391348, 179.01933225309955, 196.65346789294242, 221.17746758283343, 246.7188452769877, 262.05768668311663, NaN, NaN, 91.68188232435318, 90.63940336162965, 90.61590144981874, 90.58271494621621, 91.5791290454998, 99.3015372655312, 98.83035612078581, 105.53932490891776, 123.0315936764103, 132.0029088151351, 141.01612719047614, 152.85719919047395, 164.7555919107138, 172.80919849102395, 184.79377893561264, 214.37995499118813, 240.35022050449425, 258.47633889199784, NaN, NaN, 94.36222802482543, 92.36424135825266, 92.1215902995751, 92.30682028153893, 92.49399972517584, 96.49572474650535, 100.96049469167042, 117.0661687910247, 130.94551393669008, 140.88561145754085, 155.71755354163315, 167.488397515448, 171.752934758517, 175.07053789641682, 181.16656400976484, 196.08946961992112, 214.46581797365644, 238.66797860189845, 254.22560252704724, 260.5474724198493, 266.09460468141594, NaN, NaN, 96.47330898293868, 93.88534518982381, 93.34610762657567, 93.31121073670101, 93.27315567358717, 95.04576290186635, 98.71458310608652, 111.83718673375013, 135.51181126764763, 162.20125397456437, 177.57897055814217, 208.20848464416537, 238.964029333362, 253.6235672276911, 263.7001451232712, NaN, NaN, 95.77938503810753, 93.96180594162901, 93.67939987174533, 93.64529476241324, 93.86857762717811, 96.51946807320819, 108.08182901802819, 136.43009291614806, 162.56892283370223, 173.76786434836484, 190.97256868438728, 220.5005838839426, 241.63212896906418, 246.84298553897776, 257.93866576998033, NaN, NaN, 106.53320252271637, 95.72070878269695, 93.9344895079227, 93.67699346897872, 93.87788919134815, 95.93168141531258, 103.84343479212937, 129.21042766087302, 145.53009318636276, 154.83017571200202, 169.82122020787412, 194.61902414328358, 221.68976291454734, 237.11422221644645, 251.27922630973353, NaN, NaN, 106.84799053528741, 95.66947517746725, 94.18014449621323, 93.85606158397889, 94.12165226441364, 93.79890857566203, 98.54447596882508, 98.85871538567903, 111.75895794451195, 146.22861412621327, 168.8302923668851, 195.29361390916768, 216.24897547352657, 230.91592578866462, 244.71025206113393, NaN, NaN, 106.16142380813686, 95.86512266265744, 94.55576984162941, 94.26365084689394, 93.97370119273862, 96.02807778590467, 100.69929291826809, 101.9725250647333, 114.29352582248869, 145.47397740452445, 161.25613868630563, 178.02604090797902, 197.47982715572172, 209.11067064694103, 225.80179914330392, 238.26949229598372, NaN, NaN, 104.15806082764693, 95.3271259302749, 94.12671935175946, 94.09528787874613, 94.95391628423303, 99.39183904467318, 97.04386968711302, 97.03503951055059, 102.3076651258533, 138.53656374122852, 158.0031639334594, 165.75345510733953, 181.58710803060205, 198.7610326492349, 218.05476561120395, 235.27592050888805, 245.09064760219567, NaN, NaN, 104.24457559721306, 94.97262989796522, 93.92001938847817, 93.88951728387059, 94.89633611964477, 97.24310669435089, 96.98099997920148, 101.07623883155712, 111.08889356649824, 140.98866166308343, 158.53024636172424, 166.06885321830308, 189.84410121655748, 217.8755332430163, 240.01760066928395, NaN, NaN, 103.70655141003537, 95.09853009604291, 94.19775485847444, 95.50528175781348, 98.15493735909273, 97.93260890139543, 98.36460569511443, 102.32316542662802, 107.8124968211687, 133.20061793027125, 156.23682348850272, 164.24601324326196, 188.8154814805142, 215.12417162165187, 233.46557536929063, 247.79252692683696, NaN, NaN, 104.85511347509772, 95.36458758621828, 94.24275400433478, 95.10127675088003, 97.53810084412356, 98.19112000376086, 106.11893144813638, 133.05904334992383, 158.28285202270098, 169.06006305221163, 193.19162308041254, 218.98019940332784, 229.88339161153868, 253.91293159804508, NaN, NaN, 101.87656661160764, 94.59091761199645, 93.57954387941915, 90.92361823019944, 93.5490937385409, 96.50993835879872, 107.0755128609435, 129.5597959249395, 154.42845839671074, 167.44939981102618, 173.31332680093416, 202.7414119471723, 241.9876489055798, 262.03680963442275, NaN, NaN, 98.89330727285018, 91.90523683732589, 90.78262456781316, 90.38723555092486, 93.1248434590008, 96.41376674659153, 108.72380857197925, 122.84363390059485, 140.87819999199976, 160.2138370799741, 169.82908588040738, 180.54919903420813, 196.07593531062602, 217.30126091568792, 238.70224825374055, 257.35476196907365, NaN, NaN, 97.04078614991998, 90.74144294775486, 90.05969907835384, 92.68565400413736, 94.31905093685293, 91.66269193620147, 109.8380926000999, 146.96414068467556, 170.9025930788316, 188.0302395261078, 205.54397386669095, 224.3054373847348, 252.7747242529244, 266.72962795531464, NaN, NaN, 100.78236363552347, 92.24348641565568, 91.63568610808049, 93.07740386308556, 94.8232334451181, 93.34273676064491, 104.78369634931423, 138.64991734945932, 165.78124897014646, 178.23226163607217, 201.662969073541, 228.4546157898716, 251.03458361187768, 267.95179562341315, NaN, NaN, 100.15321236714075, 96.02373515055248, 97.03339422389253, 97.25920522397325, 95.17177217706183, 103.39328695176035, 118.56490673607148, 136.3217006229665, 161.6475404353451, 178.23262478300808, 188.1440321377364, 218.02814233781777, 243.52229152244095, 266.42637840166765, NaN, NaN, 99.20706984921651, 96.25558994844498, 96.23528173525402, 96.21273830490966, 96.47822369445944, 96.18863083114705, 104.11536833929095, 113.22818848175436, 149.16046498151735, 168.0482291903022, 182.03555216520982, 199.64995017673087, 230.13055858893597, 257.83243969750424, 270.84147479871933, NaN, NaN, 103.71755200443555, 98.99991230161592, 98.68375572261284, 98.64954480471194, 97.15701235460118, 95.40021364940662, 110.9791435151389, 137.43939673688422, 157.76727461451188, 168.99602297989978, 183.92425791592726, 217.1105809184295, 254.40156309312957, 270.6649301431792, NaN, NaN, 109.37010600328163, 100.76061861520886, 99.63618843366244, 99.60754526506142, 98.49510995733218, 101.153775200827, 114.82172197792319, 126.95194197313447, 145.5262371792748, 159.8794543051812, 174.97105137013412, 194.42062448299595, 217.25376963535646, 244.14719799422153, 268.0035604548532, NaN, NaN, 110.11820479979231, 100.99244363396375, 99.50575025640036, 98.8988066094904, 97.12628739780303, 96.82344188715165, 97.098645874968, 115.62456301762202, 141.54297845209507, 167.55911215870697, 188.90338334269165, 218.75278235548456, 253.98747020363123, 270.59192355301786, NaN, NaN, 110.0690044180436, 101.05673116284393, 98.9921770818486, 95.90414904451465, 95.88354191695255, 98.69815885933161, 119.54883076424746, 144.82155211325474, 174.0676284228883, 195.66816390711793, 225.41336665768983, 250.69006269190973, 270.97688301420044, 278.04758444264223, NaN, NaN, 103.64939995026607, 99.01305488984389, 95.4215564900848, 95.66217673211655, 96.41478495314333, 99.49112238929575, 112.86578473007582, 133.74647024207587, 162.41927452787687, 183.66104455293177, 192.43873619896135, 212.87387028659847, 235.55720760517497, 261.8970107172451, NaN, NaN, 106.013218943303, 96.01658833291597, 95.41641237995024, 96.27737962090545, 97.43326057050804, 98.31577565694293, 101.8339253863028, 117.99912698719986, 147.72704394168048, 180.3463464158773, 208.91361549310722, 243.22735874443612, 267.59378652914666, 274.69873375755856, 276.18204473710205, NaN, NaN, 98.9703584340724, 96.39022181276887, 95.64823345227062, 91.95277452320843, 90.82065220975308, 96.6834106489166, 114.3451660300404, 143.75816277984373, 172.59534764053933, 206.84334576906272, 249.7141270499443, 265.7787518559245, NaN, NaN, 97.81687825336222, 89.86967163767422, 89.25981763728196, 90.41344600375041, 91.85700954382749, 97.13275152817542, 106.83800510690988, 133.60857999279855, 166.6751518192816, 202.70745860585575, 230.40560427327267, 260.1829715169543, 272.0254773438911, 277.0653991911708, NaN, NaN, 99.07010692423005, 92.45817398989392, 91.70561212006912, 94.61402432187543, 97.52994516449147, 99.34884477042435, 112.58284111571042, 145.32295331764854, 174.50157652101666, 205.80743438194375, 249.80897368034672, 274.30428155064345, NaN, NaN, 93.67108545061069, 92.34587336931459, 92.55467544504315, 94.2953039951763, 97.3672958069592, 97.56892031623069, 97.77693679703822, 103.9445440878197, 118.94471987703417, 144.76230464774443, 169.95249830198404, 190.24593403395997, 213.09364856324893, 240.604623256144, 257.7791050875272, NaN, NaN, 94.55281930435908, 95.52986776368773, 96.8372640499053, 96.48226311707764, 95.13288151703183, 98.09713723826266, 122.25717309448758, 158.03144011915776, 183.020165071868, 221.99725027934173, 263.91521812885816, NaN, NaN, 94.2707118714562, 94.62305498688522, 97.1787462657961, 96.4194949460783, 94.92646802545974, 97.11080407379582, 100.40559597978083, 120.62339542044447, 150.0664583903897, 180.4462280999212, 224.8187632948024, 263.136848931425, 277.57192551459826, 280.15068414882194, NaN, NaN, 94.15901914982234, 93.70478089909379, 96.33216994031214, 97.18563717588012, 98.0426803694603, 99.33663949433661, 104.62522497611613, 136.434022839897, 174.55953617325605, 226.870171926726, 268.0036126946029, NaN, NaN, 98.96064457217912, 97.28997712820382, 97.6020986608493, 97.24369531838794, 98.54668197505745, 110.44034117128562, 126.33693234066897, 149.5581447136665, 177.1753845385794, 214.09592014477306, 253.60588419195776, 274.6996819633409, 281.1017039703092, NaN, NaN, 91.93807214998274, 90.64127590753053, 95.7675030552042, 97.28089967174168, 95.19873451846273, 96.47421959238306, 112.67271964212242, 135.6241159342426, 163.50925870570157, 194.98215072780803, 217.93116360970035, 249.7429039245426, 272.96861309209834, NaN, NaN, 96.31163324386962, 93.31818865914825, 93.63041333534804, 95.26213467660159, 95.55962853423684, 93.22531960284319, 99.84985614140078, 141.28967442983156, 174.5135805925492, 198.9161285889819, 218.73010137780608, 248.57968378961684, 273.0364057021467, 277.43929060178215, NaN, NaN, 95.20107298519821, 92.61446814625829, 91.49002772508666, 90.36000676910083, 89.6021226337471, 89.95032888403593, 90.66890332700329, 116.80156018418712, 159.89526219111386, 192.55984827614063, 224.29956639601687, 261.5115580600842, 275.9675146185925, NaN, NaN, 97.80808266708075, 95.21669071817337, 94.46094832963544, 93.32731023336608, 92.19973350407818, 91.83012512195597, 103.58721533522888, 122.71538842843954, 149.26444189530028, 187.15740662185013, 230.47432953046012, 254.15754349462296, 269.36592467949396, 280.4931921513286, 281.9489605079449, NaN, NaN, 100.16816295708023, 94.28241983565908, 92.79467800427342, 95.70486166840398, 114.44892346297588, 132.87077121239338, 145.04558438727722, 164.91186956344148, 180.39257767812464, 189.26430201339963, 213.99407198706, 260.6809879366423, NaN, NaN, 99.37990065014513, 96.78892178566173, 96.03788486844213, 94.54244748871126, 93.78314605844892, 93.3865078393137, 103.64723505428651, 127.1974166052477, 153.36102467657756, 174.36836564382298, 183.98700232701952, 198.64971704018302, 244.61985201740805, 271.0028339844235, NaN, NaN, 101.574652365273, 98.03377395379621, 97.71452253499764, 97.39213581685577, 95.89813991610878, 94.11053027627548, 95.2863487388184, 108.49913250400708, 130.60356006759355, 158.02627299140224, 178.09295404035814, 186.999970385412, 204.42993572509337, 240.92041221566808, 273.6119040830309, NaN, NaN, 104.87737911814196, 98.17536827811138, 96.86937027569405, 94.01607364744089, 92.96788333045247, 95.27153473395488, 112.50654862562439, 141.38171329329842, 166.9309520963917, 181.97419836035476, 196.5984809484298, 211.79024193706402, 232.43557064068025, 260.0143986380966, 274.9422096083315, NaN, NaN, 93.08996650819118, 93.3742536710516, 93.94246946762075, 94.79538279596564, 94.76643755179111, 94.14898668319799, 104.16477688602677, 127.39200819845034, 150.6569449517056, 170.74224465057713, 188.3777029575889, 216.7695026124303, 251.37926406439902, 275.8509907108536, NaN, NaN, 93.12406073603876, 90.9217120094756, 91.27431852393795, 92.35534863665625, 93.43250682581575, 93.77179670505053, 103.71158294057891, 119.88111151919777, 138.98620529544849, 155.92114453793914, 168.487060573843, 181.06303643115842, 196.8014329905639, 240.86292441149013, NaN, NaN, 97.34828896953609, 93.29880306740667, 92.19297730908924, 95.10565410901854, 100.2324794883717, 97.65642701396048, 107.22923387994084, 122.31744171385152, 145.87432352485905, 159.13568165578573, 171.35803088125402, 180.62141277788834, 189.6264075600786, 225.46028210167842, 268.3425865133572, NaN, NaN, 98.02905435844933, 92.43536839980162, 91.24440390288211, 92.98467605091678, 101.52558035305881, 106.247057440456, 109.47527779882137, 115.03468757882172, 130.3283000764562, 149.75964708850148, 164.8403896586005, 176.14409054673996, 194.64630316392547, 230.79280766754252, 264.77583052334836, NaN, NaN, 95.06988008697925, 93.73146969711331, 93.48747576412869, 93.67881907026907, 109.76383481539294, 112.4583561828094, 105.21037824365627, 113.14956203188765, 133.03006940242918, 156.7141078957011, 165.63580065096795, 172.6396795259118, 198.93416592448938, 214.9243147304285, 229.397791555803, 249.06622621953218, 265.0154369596538, NaN, NaN, 100.29782489736971, 95.14199689996101, 94.34686993437671, 98.68604198668713, 116.17288427121633, 122.60595254693693, 129.04989430107668, 124.737201089631, 135.54969936136538, 151.03829727094225, 160.89582484904128, 164.07422711048645, 177.12666330928892, 204.81395885694985, 234.01477053470538, 248.05878931507073, 256.342344061016, NaN, NaN, 103.60443748019446, 98.1913272979699, 101.24744155512002, 122.82167321098962, 131.56606673527017, 132.0829464106178, 138.25956816502008, 147.03189981411592, 153.55593153275947, 158.510463164328, 166.0932018264849, 183.9171995702611, 212.0446662366661, 241.41304400239483, 256.32285511682215, 260.7747379961987, NaN, NaN, 106.3510936253345, 104.56724205146283, 104.98374280715049, 116.2137061629585, 121.75453295446306, 123.5075952669121, 126.81850660803609, 130.7681493410174, 142.475543880572, 159.76483455394268, 163.1112807918516, 173.37397235337932, 199.1676593445456, 225.29173007018065, 238.5338579103937, 255.23973731652313, NaN, NaN, 109.94126103803211, 109.55478512456652, 114.87040449607689, 118.38594130523866, 121.69177136985604, 126.85304477153628, 131.6136869647961, 135.66028696284337, 155.7444795973521, 168.6961050227704, 185.548746155964, 206.09880826395613, 220.81789258880343, 234.07851740794246, 246.8549078673989, 256.6071102624342, NaN, NaN, 111.30370811185016, 109.99871505198077, 110.33903325911552, 112.35605135435492, 115.67855710505336, 121.76197348789107, 128.38906501534183, 133.18548592772024, 140.73374113479767, 158.0266246130809, 174.32179381159287, 189.29954905852233, 209.49354570120374, 221.1532956697316, 231.5360728006491, 241.33086197146488, 253.40897940806286, NaN, NaN, 112.79977660972395, 111.01693163387169, 110.99316958883271, 112.08087356348794, 114.5358767308005, 120.28586516205425, 128.47070560624687, 132.86152482592877, 136.18020901503735, 143.49558842671658, 167.43862287380867, 192.9347951827229, 220.18239612583827, 236.2014033254948, 243.33656524112737, 250.17390215787808, 257.07564670030945, NaN, NaN, 112.13864112854253, 111.35624538553125, 111.87059776268947, 113.41787934805157, 118.5952142235708, 126.34135337766351, 130.71112650208525, 134.03649898660913, 137.90282895965936, 143.5750314188364, 149.74524908019907, 160.5834624284375, 182.3496196876234, 213.80038895194474, 234.27358334065715, 244.0182210269681, 256.8817439776033, NaN, NaN, 110.94856209770465, 109.90072023210612, 109.87417458516106, 113.47743917760188, 115.55228718284309, 119.16660656529106, 120.18313949317289, 126.87696716147238, 131.50609346888615, 134.58201447213713, 137.9097584582417, 142.2858657023255, 157.28118328057883, 185.54284327244108, 218.06269110787312, 236.69734677749506, 244.54467135633516, 250.10633986616523, 257.40033407779026, NaN, NaN, 111.67940839599034, 110.55875627356627, 116.71609702259178, 123.06507343070471, 127.43768814578601, 123.47683466889768, 118.4449533217564, 120.42129473867918, 126.16783788258132, 131.90275242972587, 145.17499561261633, 158.45076937663464, 176.28136558315174, 202.48207765485847, 224.55234946399344, 235.88209495113603, 242.83039070006285, 252.29576095248402, 259.8272777092664, NaN, NaN, 113.00303035671709, 113.72088026202472, 122.93272348699303, 122.05445798105656, 120.04513577718525, 125.40087434162477, 133.13159609416562, 140.6652576280664, 162.53665463542578, 175.6975083011513, 181.48225326410528, 191.46683736593434, 207.9610244850971, 228.80132329986117, 240.9904125710269, 248.9092787542927, 259.11805991907994, 265.11715097624614, NaN, NaN, 111.32887913185232, 110.93974614608234, 111.46301085899223, 118.42551152822384, 124.51179396240953, 121.56740024565532, 120.28611260847792, 122.67301612829182, 129.67626150488556, 137.23844139747143, 154.9390765567971, 174.40010525622543, 190.69866658762209, 210.92660276316232, 229.74620882399404, 238.39815294016975, 245.47109893507871, 251.51007644984506, 260.7166336052065, 265.4433773790822, NaN, NaN, 106.47579988834548, 105.36248704167416, 105.89806837142064, 107.34150888810447, 113.57640612784915, 121.89175786971838, 122.0933011317277, 122.64317449628406, 123.35605881103452, 127.43523489762828, 138.6787804294074, 145.30357093100992, 166.86589047538703, 175.05551902558966, 191.237362833394, 206.41806665210007, 225.32797843331156, 234.56053735300767, 241.00720744896356, 247.29496746796724, 259.7686010551335, 267.8633258203083, 268.26268304865243, NaN, NaN, 108.1606426638745, 106.31679680267358, 106.48206823506035, 108.68573880500183, 115.11582656877377, 123.21463305860371, 122.4892934443523, 120.8290362280541, 123.77147571877194, 125.61071886924235, 133.00763437994627, 143.72278149436005, 165.69614136098517, 174.04405239927522, 186.62163904922593, 207.22423938873365, 230.16425706678794, 239.760504682441, 248.7088786016208, 256.91809237593293, 266.2867957675284, 268.43963298172923, NaN, NaN, 107.03142501399387, 106.15223050316844, 106.38356762614069, 107.93659560504476, 112.77185506298538, 122.47000430979485, 124.89556538321274, 121.83739266978475, 122.9485582632682, 125.14903874825734, 129.32465731995782, 132.4482021931286, 137.74069173289385, 159.16056208407431, 171.4472454985728, 185.4432070684014, 208.85219435620493, 231.94899040708887, 243.11581841286733, 251.0046136665481, 258.84420967795756, 268.5083126972599, 271.062055780267, NaN, NaN, 107.18847685748737, 106.0210679650526, 105.44820627510195, 108.38862671509308, 107.79891321872526, 112.495362452325, 121.59252320779751, 125.6983944074407, 125.08830175061843, 121.87557477623989, 123.06002401768062, 127.75919270283394, 125.45948385904975, 127.20236803798953, 146.9201125194213, 167.96313864687275, 192.06568536292042, 227.86728063208633, 242.3649554450183, 252.39721581303687, 259.97290220079, 266.2091175103642, 270.195534753067, 271.3098768099678, NaN, NaN, 105.78586859845993, 104.50654057713919, 108.62970212307278, 108.15586515162556, 106.34550211184018, 102.4927836469974, 109.66994493708897, 122.26172048628547, 123.81435239535239, 122.5059752894127, 125.32714332015125, 127.38254484926293, 127.17553629081735, 136.71458417113055, 156.28630133125716, 169.5070364099752, 180.20104691653742, 209.58266872526397, 234.48646884255083, 244.85792505709546, 253.34959576045924, 261.08369526472563, 270.71305807304446, 271.9141210232608, 272.1803136303111, NaN, NaN, 102.8475487901395, 103.39468593909321, 104.68643746790937, 111.67422786522775, 110.0181130741554, 105.22924732445011, 101.39504358962034, 100.65047352141464, 109.61897720364905, 121.5662922511621, 126.18565425521844, 129.5098784830033, 131.75364726536736, 138.19791941383755, 160.11617235813807, 174.62596557029892, 190.74466126942306, 213.69614620180812, 233.1356388735677, 242.34507569606154, 250.60527772636732, 258.47047952327557, 269.61846154769887, 271.805742056873, NaN, NaN, 101.69310573365999, 101.09943099247623, 103.4347368497324, 104.57380192138396, 103.98117716082203, 106.9016299589511, 108.39156467030541, 108.72233677572885, 105.80401210262963, 113.11961940563023, 120.14850881238532, 123.11707211474145, 127.54878119677808, 130.2487818439919, 141.47300969401263, 161.80052155151134, 171.606088294757, 187.67581859208588, 220.9518531240448, 236.6449950267769, 245.6366167139833, 252.3224988356177, 259.9178745661306, 269.06236002383514, 271.65160428608203, 272.0524826099405, NaN, NaN, 96.37354082920963, 97.64800725761306, 98.72914040663088, 99.25468868232744, 100.33557369152506, 102.36818949957103, 105.3200620586793, 105.35166992182097, 105.18766355531639, 107.77129774233565, 118.04034823333815, 122.45426860714953, 123.22094138614949, 128.590213657902, 137.07083649886545, 142.25654032678065, 156.6584959033157, 171.0628155526644, 176.32236805153696, 195.0575999560118, 221.53639965552713, 237.2632239396052, 244.01336784719706, 250.3070464858259, 256.3381854022164, 266.88525206253564, 270.38524438912737, 270.9406092653689, 271.19109504191346, NaN, NaN, 85.6080377664338, 86.25644109557238, 88.55438676563391, 93.71965826170172, 96.68613798329169, 98.31374796515061, 98.84317756494045, 100.8266846146723, 104.36821539102905, 103.97844807750133, 105.29779055517616, 105.28741830781252, 111.20968576061009, 121.20440729697947, 127.83014719620618, 124.54030380185692, 124.703177036974, 128.44321692525745, 132.9655031890266, 143.58220531835667, 152.01439769888543, 170.15082763262237, 182.05825875308165, 206.60773769839048, 231.99932107804224, 240.18524572764488, 245.49992822986195, 252.00341414652146, 256.6078375802348, 266.3115143793675, 269.9111363920209, 270.3119383400284, NaN, NaN, 67.19700253713133, 67.87016973097282, 69.05613798796088, 70.58389526524653, 70.99794367553483, 70.97238026715544, 70.7274675653148, 70.70363842908843, 72.15773525332027, 79.12581321769073, 81.97683795850425, 86.15423435621442, 88.40803769272149, 90.36980933358258, 92.86691631766949, 95.28960855207146, 101.39634235813702, 104.50320485190541, 103.8995691485975, 102.62472087304018, 104.80003342237495, 104.5913646164092, 117.80680207880711, 128.1879000973308, 128.9081663702448, 134.72586240318685, 140.2580438089782, 141.3482751470646, 154.84498501357643, 179.31709198837518, 195.26422765780202, 215.94678857463845, 234.66737744298604, 242.68589179246302, 248.23863248443058, 254.07846432327807, 258.65591296135784, 266.7064093024592, 270.0856566131277, 270.097434240736, 270.2711757650306, NaN, NaN, 41.02666115030212, 40.95374062966509, 44.051507086461974, 48.168574359244616, 51.32716228647058, 56.10673674573061, 60.88475768447749, 65.22037229409419, 67.41398618452821, 67.48454473698153, 65.56856528765269, 64.31142986284969, 62.39041478216428, 62.82406148564142, 61.049094171716135, 67.42855279297423, 75.64137219881115, 81.06472355225188, 80.02705228906294, 82.57588995304391, 87.03348155067091, 89.08413968600777, 91.1320900921109, 92.57977761706692, 92.00334025388771, 95.6695271970314, 103.43783859648018, 107.25574852873076, 109.46830731763066, 111.38457154690903, 105.8143844880299, 117.44165035951065, 132.7134283947078, 132.27332319518237, 126.70828311789937, 128.51833149055676, 132.24080547735682, 136.36701190319138, 141.10501256535784, 158.06675349381584, 184.7448318481749, 199.0646262007076, 214.97566801072594, 234.18840914634148, 244.6800138719717, 250.7077533827263, 257.157252915611, 266.4707271723637, 272.342812772222, 270.86898514855784, 270.46249253646477, 270.06640753736735, NaN, NaN, 23.340041363023794, 21.605483770703387, 21.601221692273054, 22.114415755450278, 22.697534984443106, 23.505764974972536, 27.310555869313433, 30.10619538451614, 30.72375218995388, 31.416077157385576, 32.88680088781618, 34.576236550255125, 36.192072573274224, 37.32401716624132, 38.97420557884014, 40.736092950082906, 43.82301176185103, 45.762193310840104, 47.11250810496838, 48.572065869231515, 50.77591460937248, 54.37081214320227, 56.341892992471074, 58.90192457208552, 61.985022743725224, 64.25061326823459, 65.48123252149716, 66.57829164074201, 67.89405519545876, 68.40019667555508, 66.56716914517028, 71.55625061564076, 69.34753619096243, 69.77493519079817, 77.32129785999852, 79.36746526410913, 79.21012389158376, 79.78001851440854, 81.6069074623295, 84.96415268918284, 89.50493788043273, 95.23181263275964, 93.27566700936903, 93.05991442595482, 98.7854074756556, 106.71129838084576, 113.97451047306792, 117.27406195345534, 111.77892391449252, 101.67753697561491, 110.49840789238976, 124.40303506752659, 126.9014950137134, 133.58682912986282, 135.80269993584548, 139.99796806407073, 154.5929916107664, 178.94401690187655, 190.6373127651319, 202.32418604921372, 228.3784710641277, 243.7658151576933, 249.89669005293976, 254.61743522624508, 258.0835272795226, 262.56490317700013, 266.68713356359626, 268.8297796107717, 268.41371232372353, 268.0146629419925, 268.13179874479863, NaN, NaN, 21.579911253560415, 20.875943556174832, 21.093648976118224, 22.681741164341265, 24.41281935871373, 25.550422124144603, 26.83521666852041, 28.41443682743474, 30.066804969346446, 32.01553645528638, 33.59130476935856, 35.099940024487054, 37.23029063834145, 38.50995062978133, 40.640410172902655, 43.09506430051629, 44.481426465791415, 48.19177602641722, 49.87459216390853, 51.296895024506526, 53.38539890135281, 55.07221902143315, 57.27047451659107, 62.18352625070704, 61.077766528825514, 59.67203185480309, 61.05916835751591, 67.87780218581537, 71.75925748343346, 71.16922781526611, 71.96877014263751, 72.70200999982707, 74.83164814660981, 76.58353186098283, 80.01313254873556, 83.37935640454558, 87.10716616094695, 94.36681058391116, 94.9418799843379, 97.13617220574825, 89.2204154824792, 88.11257509385574, 90.31853788913035, 93.84529382267162, 101.10740679123444, 112.12693644211573, 121.61186599235852, 120.96124076119509, 114.60050910272213, 117.01678315509706, 119.0179758638485, 135.3578573833212, 148.41249311445688, 145.8832856130221, 162.72049534907867, 188.9744595693303, 200.3259358486916, 218.2939682875513, 230.55217440178663, 240.8990966274492, 247.2532494664965, 251.10620482790918, 258.777560285451, 266.58474451309183, 266.21896304036767, 266.8615442535407, 267.5840234070306, 267.7205178512613, 267.6886565812068, NaN, NaN, 20.848133240481246, 20.476000247116886, 20.730357786374228, 21.574149855366393, 22.268728379305077, 23.074309903779035, 24.13774243636371, 25.4221150897081, 26.55812028930099, 27.989606530075935, 29.826346574416995, 31.88214514351334, 34.15580331541726, 36.02440255508969, 38.29962942151814, 40.98377388346037, 43.40848843985132, 44.28548339431474, 45.74797115552986, 47.17305977053023, 50.00135841261063, 53.82016894146971, 56.833896728638116, 59.39453834122882, 62.10058447137175, 63.12048978859395, 60.980429467056936, 58.62213603272767, 60.22761467586193, 61.686581409025926, 64.10840744067652, 66.1553551364043, 68.79353588227428, 73.55958489280772, 76.8567236413661, 81.76129407173417, 84.0975403578768, 83.43068119729453, 84.45274302459032, 86.06414389100838, 90.42881982524307, 98.48030653833885, 106.2652999201663, 114.64399104061903, 119.05970393290984, 137.4254004904361, 151.81226402858167, 159.46061305576868, 168.43602780237038, 177.31350965489423, 182.8599270639855, 183.37367327161368, 189.80714778831828, 195.0101202694171, 199.97629473213854, 199.3828718967688, 199.9306444606271, 199.43850690233157, 216.42232732601556, 233.6738060883673, 243.70015631660283, 248.1966731323464, 251.5078999450595, 257.45728565516754, 262.84668740778534, 266.8363241690232, 269.86696973322995, 268.396679096432, 267.62837891713497, 268.3396350003234, 268.04674212991324, 267.6046981385613, NaN, NaN, 30.06280123158788, 29.177467794224835, 28.807150845198045, 29.76013653443026, 31.818183592134098, 31.15350764392423, 31.627600201197826, 31.21845327229233, 31.10120990438445, 32.200407267077104, 33.295751897509305, 34.39105493594629, 33.98093425497252, 34.12156548436516, 35.290905955412605, 36.792554661841194, 38.47897526148468, 39.7970952157268, 41.18475837746693, 42.05667299760408, 44.921039639051784, 49.217433647595584, 55.05132014520808, 59.00570167518978, 60.21568021739969, 60.873428075905515, 62.410022935078864, 62.40471480897552, 62.6175874436829, 67.89511611887518, 70.86220805411656, 70.74065523210955, 73.48417526414285, 75.24147560414654, 77.32065810202444, 82.25954467298654, 87.31454226016257, 92.15599957013926, 98.96504456402754, 109.40214476971038, 115.14927638056683, 115.88243883644876, 118.07824262399711, 121.58013265549415, 128.9220720429345, 137.725451136089, 141.00814310426412, 152.2254923324186, 165.48339987959002, 173.2324377865777, 177.2794437436828, 180.61238654622122, 181.84133739658654, 186.95973316950924, 192.83259437624093, 199.33504971564386, 206.32348054678147, 203.02098967690847, 215.47206837478285, 236.9449759872077, 245.00200678878505, 249.0200137209321, 254.02682908961296, 260.3435515478635, 266.691900618401, 267.2867765566601, 267.5167331463734, 267.4265517442491, 265.04700175747973, 263.1342427302543, 261.9612877708938, 261.5516158232992, NaN, NaN, 22.324686471007144, 22.251447663741242, 23.060739545479873, 24.161852100117038, 24.597115046805527, 25.845730810922433, 27.683635021503637, 28.56133840473715, 30.102195400263813, 30.759888842274314, 30.238843933777424, 31.11877427920222, 32.36438424348612, 33.46065352121008, 34.55773026232876, 36.0234294924611, 38.00301493207614, 42.779214034783635, 45.638200577599086, 47.40373595935666, 48.905431972126294, 50.11350846906584, 51.98074262436004, 53.40446323634245, 55.15901740915748, 56.804927319685206, 57.89834401012087, 58.99209883137455, 60.744635512756616, 64.36924508655167, 68.10703242990972, 70.95914214990681, 74.14580417393414, 77.11187808603465, 82.27373404741678, 89.52794991653491, 94.91531520792093, 104.35881374916184, 113.9077404672191, 112.46992938110563, 111.7265748084432, 114.06443796504058, 116.10528418428278, 114.92680986287327, 120.06748192309816, 134.29177727848412, 146.0322102078369, 155.29978637630913, 160.0062717176555, 163.84798195677, 159.98619138233127, 161.1813629073043, 171.2690203905912, 182.09077881591443, 188.96573750587834, 195.06562932132408, 206.13960100068186, 210.74299571830042, 207.12620023231253, 223.91575044687386, 240.39346459785568, 247.40841449521972, 250.65380318464122, 251.83257010596185, 257.2926120811862, 263.1156144388741, 267.50017091719377, 267.73497006825363, 268.72442060526924, 266.47965120210927, 263.45106087379327, 263.2530987307489, NaN, NaN, 21.993317599769515, 21.400635181045747, 22.50343977885047, 23.67565879736388, 24.999178308694432, 26.249159513021212, 26.425748141845553, 26.9005484938352, 27.81442833116619, 29.246382888434468, 30.78757659992364, 31.958887381737647, 34.198533093205995, 37.90647041391846, 40.68953343352426, 45.05829979498612, 48.13859421488489, 48.01750246485684, 48.045596914221896, 48.58612062221048, 49.5749700435094, 50.23306109531019, 50.44363899187176, 53.40991030279778, 55.82428972196866, 55.92518000111938, 57.461391436871956, 62.520723805486945, 73.0866719949553, 86.1795300293292, 99.04073774207801, 110.0328376433314, 114.7591229936764, 113.98688913873526, 114.8643450464075, 120.24432106968067, 122.65490435145834, 124.84235241635193, 128.2316986756471, 133.81714287509462, 141.71778862703474, 143.77374774786023, 145.98412647112764, 150.83287547510182, 158.47864963384043, 161.60298161792673, 163.52382195378334, 164.19266251580052, 170.25113559367276, 177.28264724023873, 184.05303728019652, 190.24627663453745, 202.28989441959212, 214.08835734696615, 209.49867962827986, 208.6027908024011, 226.86075529727958, 243.58909192511143, 249.51287631320665, 252.31173116396164, 255.1510951566605, 259.63034357336045, 263.2662215880788, 265.42632704716107, 266.57535986690425, 267.90226263537147, 267.6951871995569, 266.3155387953393, 263.933188334947, 261.29477787455863, 261.1664481028937, NaN, NaN, 22.43757094678572, 22.841073704985156, 23.720648958709948, 24.45254295285588, 24.927219570321963, 24.994713267298756, 25.06196892718591, 25.27785285545125, 26.046250190318307, 27.1819797763098, 28.760212745308973, 30.261998258161373, 31.396852743909037, 32.60505571085816, 34.58537426771094, 37.92270210804083, 41.29987311259714, 44.26509114009679, 47.04877181084891, 47.04389174032615, 47.3726557559863, 48.286231744705766, 48.64238258700184, 51.209219707044696, 54.50974295536427, 57.07274300607169, 61.107215446960296, 65.8787431512853, 66.97383633166733, 69.35359999194434, 72.09631800634672, 77.22656137978609, 86.20445455595788, 105.09287264226958, 108.02373557802086, 105.99502243838826, 109.2793743514567, 108.53219037382262, 107.41939565989966, 109.25709402393372, 115.26338687235004, 132.5728609443224, 144.46120981683492, 146.3872996485526, 149.3352862006971, 161.2350154165713, 160.97111683195803, 160.3085207286257, 162.56965311738446, 172.35712205348003, 180.85945700689797, 187.04752196163363, 197.3398935916904, 210.3740635269468, 221.06649448891523, 226.02278991722878, 232.15901497597895, 245.69161869537103, 251.7180071673997, 254.91444823271922, 257.40022807288284, 261.4979782744288, 263.7321291992935, 266.35191250282537, 264.2467694626329, 264.7200746249849, 262.0791188268721, 260.6405583247745, 259.98212051027514, 259.9141313918188, NaN, NaN, 21.844408959722436, 20.072798929484208, 20.437887936456608, 21.243417235689602, 21.901429634990052, 23.000881458939578, 24.763423003556376, 25.71295815743443, 26.00113372432485, 26.289705030637098, 27.68337828959114, 29.294498351909315, 31.715351429198034, 33.8436269612513, 35.3088029600075, 37.214656558995, 39.12176564967688, 38.82771806734682, 39.554381204427465, 45.491931853918395, 49.15535159579706, 51.68661151678532, 53.00489646824688, 53.7710838923039, 54.20051861423753, 57.50035426164693, 60.139054845416304, 60.794075585301336, 62.99047524914639, 65.95712263662655, 69.15313274390802, 71.01485980511717, 74.19403964469574, 80.23627341473227, 87.0529533273177, 88.36195763727113, 92.42767005221646, 96.27483115694382, 107.15247805510074, 117.70427485529122, 116.20622726472452, 118.56755981696152, 120.91169480558604, 122.52587977843476, 123.55789829164097, 141.61747946415008, 158.07166845616322, 168.5269393125157, 173.66787795959183, 163.45197434685667, 168.80243064668383, 175.9566731214144, 176.65609606421245, 182.327644188133, 195.9384045976479, 209.7640348502202, 220.6752844209115, 227.44330149305284, 233.5111896733467, 235.83405716100063, 246.7408504058636, 256.40097162996886, 262.0477607750118, 266.5215527141936, 268.28594185512196, 265.61014449058615, 267.4091033788224, 271.5508796487707, 266.8503198390046, 260.0654707937879, 257.49795431197214, 256.6905024758389, 256.5246849537994, 256.26986059214033, NaN, NaN, 19.632020773908454, 19.29706499665283, 19.99467636252137, 20.615908152225742, 21.38556633423091, 22.560028594384068, 23.58747342133771, 24.32105380523108, 25.60380637939699, 26.371589591388084, 27.02919087421101, 29.122158253063883, 30.846345843226008, 31.80052351296335, 33.74448126755437, 37.15545802633252, 39.24598625979507, 40.26878084172912, 40.45161242533566, 42.943409706111716, 45.36042780388014, 48.659479030723425, 49.831141372106636, 50.26383922739085, 51.80063005746542, 54.58362300409891, 57.14651259130476, 57.802782420090345, 59.044507173762305, 60.431255558193534, 61.81830915907069, 63.57950606737866, 65.40819487174286, 67.61048858874727, 70.46551977013031, 72.73488676704629, 74.99988671468584, 77.93204435011815, 83.13806198775016, 87.08663442024093, 90.3842771039944, 93.74932025059267, 96.82257210073655, 99.7510104475222, 111.18992964322565, 118.98499696833534, 123.09506862416227, 125.44106335306867, 132.1952954421632, 135.12888929978732, 138.8089690005843, 149.10498159547592, 163.79872954092266, 172.32740060681058, 179.89748944340332, 187.09253512165077, 186.30578195997174, 189.7539755686756, 198.7449315096191, 209.09329534690264, 222.55861785335304, 232.5083223502231, 239.7709571441468, 247.72308176212417, 250.6331477713107, 254.53088336047202, 257.3642425147286, 259.14451725802815, 264.17711363035517, 269.83908443844274, 267.959951625141, 263.6764200591868, 262.88660986299334, 260.9750994310077, 254.70604951337907, 253.33917381883404, 253.29631438526607, 253.48206334163794, NaN, NaN, 20.923326399944166, 19.852008944353276, 19.850360609956255, 20.400427230640815, 21.05922915084177, 22.197260934691993, 23.001675597896384, 24.65292670871223, 26.230109759040566, 28.691608192896073, 30.7844407517636, 33.42950504254049, 34.41674322309094, 34.37846485566653, 33.860335240827574, 34.221017350069374, 35.8674637442842, 37.81280340371654, 38.583709375278914, 39.93722462066777, 42.759496667697974, 43.78301344544867, 44.0762535300828, 47.230419540585224, 50.8213941669903, 57.27913028980259, 58.66600255539167, 63.501759514496655, 66.50603771586198, 70.31373950873417, 73.9023598001914, 73.97070825375485, 75.50719173129535, 74.10145036392377, 74.59868499531451, 76.0538239009228, 77.14739908473383, 79.1197642271001, 82.34617376764876, 86.67556027682222, 95.86793882041064, 101.43899491532048, 111.99564212420741, 117.72106623687502, 120.6802204348842, 123.78752103825303, 132.43566776342294, 140.37354979398174, 154.64615432492081, 168.94386505228982, 179.18104539672692, 185.6162062559004, 189.1254288981891, 196.94964086016748, 203.38143118083246, 211.06218375776135, 218.5951509324478, 226.12966818267662, 233.10268287620246, 237.0653072721412, 239.183507399325, 244.11512151425606, 249.41967646377014, 253.5696568401302, 262.2441924855909, 264.27647394108396, 266.99563080823776, 270.5441207501252, 267.43012690929714, 264.6446103373423, 263.265459540243, 260.18070565698815, 252.6878514008954, 251.58733688833132, 251.68839803759346, 251.73434196168, NaN, NaN, 27.456045193372642, 24.095605825353747, 24.12733247693993, 25.117009123465497, 26.438995206507926, 27.134644410340496, 29.375485808926268, 30.953957068819776, 29.700323628830972, 29.25590875988432, 29.43505124047177, 30.643433403448608, 34.42726670321226, 38.13728075588601, 39.7137280722982, 38.86200474453329, 35.95300771708001, 36.754296691751875, 38.99026311535528, 40.311176435777796, 41.664920868189775, 44.74318958681746, 48.18808624816777, 53.61991779547065, 61.6894688537485, 67.48603343436352, 66.15898475566418, 66.81830579639237, 64.45799971069796, 69.00823643014924, 75.02347990710356, 79.127232693221, 83.01335449915676, 84.68896278428875, 87.9784266923047, 94.35174371797223, 102.86204212664003, 108.06232894263894, 113.48469318774181, 116.71764038073411, 119.8651242566197, 126.0272653889317, 133.2232052023087, 140.42547547188477, 150.2701113645328, 165.13169179869558, 172.95032314801688, 180.82483330406507, 186.37953161857402, 192.53973933704825, 198.202473223784, 204.3887130449291, 211.27338087988204, 219.37689407736556, 227.41084631155206, 233.63813328164167, 239.22451245956756, 242.64095053140682, 249.48817365628324, 256.42258928034414, 260.08341753623074, 264.88635397726426, 268.18755953075095, 270.4633744595898, 271.39138310177987, 267.39906749158274, 263.46154285441196, 261.597185566326, 253.75595516144114, 250.8735383535409, 250.6843946566508, 251.02711448251446, NaN, NaN, 28.927399837068645, 26.085424486444126, 25.822871257863298, 24.824741864486484, 25.481974934943104, 25.84539991573507, 26.42972799083608, 26.864729559295643, 27.080782290744636, 27.481016308416276, 27.955479819127667, 29.423199242362024, 31.07360607787783, 31.21570293683059, 31.614238181130244, 32.343671367960575, 36.269412669593834, 39.497792226295005, 43.45935342412572, 45.43591137954023, 47.963317819401674, 52.509872440643264, 57.94119668754814, 60.87358426975636, 63.21887359797561, 64.97567869273765, 63.6560175305583, 63.9394962764098, 66.72461385427064, 67.00642702542338, 70.66787007848747, 74.76789296295404, 80.92299249718633, 86.0450573879851, 92.50168275970867, 105.56132900072984, 122.72121085639387, 124.78494544683305, 118.4728749362505, 121.55793591633088, 123.5650921379573, 124.49118911732319, 128.16540348222895, 133.12885632711857, 144.17473616121802, 164.20881987418042, 174.54822839353986, 180.6895153043182, 190.84084413112768, 198.1442071714279, 209.28806233686396, 216.46619900905455, 223.0344216716056, 227.7935143642375, 231.62498746995252, 237.00344781243274, 243.06703948666055, 248.2949601108891, 254.85447256008695, 263.01597727037864, 266.9874405194908, 268.0340506121682, 270.6031818848456, 270.997928825884, 267.5357338425868, 262.4459056837476, 260.7031972515935, 261.4577743871339, 258.6926694730158, 250.748492840012, 249.81078786885047, 250.00042557270024, NaN, NaN, 23.213624640752887, 23.799192027695575, 24.53367399951073, 23.940090151124245, 23.458414723394007, 22.830621903325763, 23.345564881778103, 24.665094077699777, 26.574167499265272, 29.145323801740847, 33.479665690547925, 34.13722577754153, 35.81828379632538, 39.52480796360027, 41.3586917726339, 42.34562698430623, 44.359798577799815, 47.47386400303597, 51.14207563128092, 51.65116443207257, 56.45411229663906, 59.60932850265987, 60.55359212308727, 61.0610748430379, 63.91990792822078, 63.02715385216706, 65.14854408066249, 66.09675479468541, 70.49637181866487, 75.76964853460896, 79.13553891678184, 83.23828315026023, 89.31842419609333, 97.15900738722128, 100.44720614137195, 103.07466771825514, 106.65978924954875, 113.47504101732238, 118.60187404313007, 120.94625478562864, 118.47853110554469, 121.58263002229309, 126.57643004995273, 132.6068441032059, 143.6463539999849, 161.01870431438064, 171.76629019747813, 179.6563121923657, 186.6481133789001, 191.546109411203, 195.31592877706538, 203.4860569828319, 212.3936616454533, 221.17125055683857, 227.82190707252715, 234.4107778151661, 240.68821074212826, 245.2911283204854, 249.75246516929846, 258.4658578692022, 263.4617334939361, 267.3935957361909, 267.9521818791791, 265.5632461763235, 264.42195554156933, 261.29481447672885, 260.50747360847464, 261.4148104055305, 254.3742072915656, 250.06269599206837, 250.07787485413638, 250.19584475583756, NaN, NaN, 36.04036047753044, 23.980277668460346, 22.3174317881965, 21.651878793566503, 20.875225675606686, 22.30610860621462, 24.179630006324775, 25.832098074292425, 26.491206026001873, 27.48111424684262, 32.00151305047033, 34.42402280071753, 36.29517363289551, 38.05443701855782, 39.70366032530738, 41.23952257987566, 44.54024686302953, 46.301967066131525, 46.18751360166387, 49.04649798140379, 51.16998309086238, 51.60417615618812, 51.817154909693514, 56.216171920622465, 58.41525474613982, 63.25507389922699, 65.1175677513668, 66.76042813796448, 69.06724628917604, 72.47446067798144, 78.7436802479462, 89.52611475576036, 95.36074601437636, 98.43474774263126, 101.95223579618046, 104.03363552612649, 108.65351668253362, 117.45124611203147, 124.60770927437763, 120.75531559659981, 120.18160984446429, 121.21413308500817, 127.22866129352546, 133.6885619498934, 139.57876003212738, 146.80868120672358, 161.70422985595636, 173.94949331365666, 181.12722849914826, 190.91788757843725, 196.02397337922824, 203.72435364526422, 214.02565249913297, 222.33584133241254, 227.5998295307403, 231.99092000839937, 235.824541220739, 242.40951480588691, 248.97677222477378, 254.55776898089192, 259.9927230029521, 263.32017455521736, 266.2743307265172, 266.20183289754624, 262.95234354594146, 262.7436451759098, 265.8438567448232, 268.1086726140178, 265.7166509188058, 262.5806008832948, 256.32303349045594, 250.52182075237144, 250.1668344746224, 250.42132656096547, NaN, NaN, 23.35900665388059, 23.024105977833052, 22.87444811447883, 23.60513968785957, 23.273231607193342, 23.638608862030313, 25.07285865517124, 28.822257547612768, 30.06978572441865, 31.246274759120542, 32.858442725186265, 35.50220105829117, 37.88960806759084, 38.91776087833589, 38.94824800083733, 41.00133932889454, 43.56947871448696, 45.66052983558089, 49.29318789789128, 52.33926543055759, 54.3152416814984, 57.83559207331265, 57.538290769243, 58.412906633510225, 61.78435793739545, 63.683023655912855, 64.5637608209441, 65.29328601751821, 66.4579407450504, 69.24076200124993, 70.2706418670367, 75.98972017498589, 82.29295153978161, 88.15666424063363, 88.59669911694566, 89.76352762069251, 93.13272243390418, 105.1660913686286, 120.4327778613074, 129.3919296298442, 121.97088054863612, 118.11873906035744, 119.44929224601321, 124.98556389282194, 137.24234544894884, 147.50510051753497, 150.06904627747483, 154.62533217012103, 166.34704643554787, 178.32330720460902, 192.39047529751343, 202.1551712819783, 208.57754893288535, 215.3897311513106, 224.6441509915523, 230.83659966851965, 235.29665536694563, 238.9946631604616, 244.54992573096465, 250.95613566423128, 259.1890651891891, 263.09769740396933, 266.25853406543376, 263.3591100075416, 260.40146006606193, 260.0377093492976, 261.5928915500223, 264.0334005417548, 266.7963217092053, 264.2905293178736, 253.55408851095137, 249.8592719782244, 249.81306993256968, 249.90284383020364, NaN, NaN, 22.621038402872355, 22.839992762098056, 22.802231347192983, 23.64462852020376, 23.864241684798, 24.340461041101097, 26.51161706348986, 28.310248483779052, 29.29923285652618, 31.096317921002, 31.940516955654285, 35.24696304201117, 37.19138504121027, 38.21649589340454, 40.49167826190741, 43.576059243200994, 43.977140712706706, 47.27729647798066, 48.079465795074555, 47.8510841376666, 48.06339140173861, 50.03847414075107, 50.91284634935471, 51.12667489749322, 53.434435086423264, 55.19415280422616, 56.84098515180764, 58.04592502482535, 59.253299834855625, 61.781349624672934, 63.31171951509814, 65.06707472420234, 67.14909995540553, 70.00281116953626, 72.63767638081525, 76.26353167808205, 79.67076990581879, 87.2587500165396, 98.47071739192208, 105.29779702646239, 104.90734273993495, 117.46664731150211, 120.36001725411735, 124.11486109759554, 129.41029068259996, 138.2575663013522, 148.87861870843622, 151.96233039311136, 147.64520292185912, 148.39213346994993, 161.29323797500479, 175.48835187642726, 202.16174466201704, 216.31737551700454, 226.32556168029424, 234.3394451706873, 242.46801826790903, 248.31859394046828, 251.37342002244827, 259.7900310610294, 263.79191470010005, 262.2234338588287, 260.4766496839675, 259.7661402627202, 259.3435386729754, 258.364660484412, 259.6771326486541, 263.8358640065828, 258.3997736097321, 249.9591225807463, 249.53555067299084, NaN, NaN, 23.399958394700597, 21.70183791226842, 21.440454526743878, 23.314755433600862, 24.27063710227684, 26.441460706271073, 26.363320073616947, 28.97278120316183, 31.251705688420117, 33.45515751554895, 34.84761963555048, 37.860254476197156, 38.84780224233253, 40.606104672846065, 41.95887528089956, 43.72192738035634, 43.75031153397933, 44.13531008915393, 45.34488920859273, 47.87589250120661, 49.118409407403114, 49.92053543024592, 51.535004397556925, 53.03334040357978, 55.41650576411234, 57.35644747117026, 59.58772923555296, 63.977457947099474, 63.391558388681695, 63.1977720547767, 66.30651672882475, 68.06215200644864, 70.44308680257045, 72.85989478690944, 76.52310244018864, 80.6636923565532, 83.03755790809791, 85.24175811332739, 88.17065110775901, 92.207774076179, 96.16646489764885, 101.16835147601148, 109.8408058632811, 119.98625754890351, 126.76076318073457, 132.70536863759185, 142.61419509993593, 149.73619606402067, 154.17629463885967, 166.9288159185585, 179.1410751762037, 195.7278373313394, 214.34614669990924, 224.15878886978365, 231.84647884379845, 237.72447879811097, 246.00780129221533, 249.45099845218016, 254.67447261219615, 263.2127136988328, 264.2890339078929, 260.8361021297084, 260.1131566958664, 259.5155184168638, 258.3452543053082, 257.3032876767981, 260.838323705074, 260.66723152995576, 251.2234562471724, 249.37408019741164, 249.4461785555847, NaN, NaN, 21.81613478015458, 21.518346633299984, 22.990164021613065, 25.15934105027158, 24.897840325644555, 23.860777156460937, 25.5469879801272, 28.634352440625364, 31.35571747711969, 33.04643024541343, 33.48530434967266, 34.95364535115376, 35.94105353608378, 36.00763196860824, 37.433461426577686, 38.74794524401071, 40.580665506409446, 43.73352438072497, 45.271870753621734, 46.29697154173132, 47.57721604104555, 49.480521772211176, 51.383012858574624, 51.82108939620426, 54.31423720870336, 57.614773190122655, 61.13625479254426, 62.45224303501816, 61.49713680876863, 63.771848187046466, 67.36935934358084, 71.62590107244566, 77.41769795281303, 82.92076365126428, 84.59543142597533, 92.72162484758489, 100.86467587195546, 100.50826099400034, 95.15678607083322, 97.41816277915905, 106.37035733997882, 106.39874696456992, 106.93259139819045, 108.53964070997517, 110.20597291242784, 113.36415633644147, 115.87900549810095, 117.11329531939873, 117.08039566776822, 117.85756899316517, 117.72877683415956, 116.64297201403006, 116.36176515545807, 116.06708390989732, 183.3086447672315, 235.50302736014558, 247.93339548117973, 253.66646881569102, 260.59377593098935, 265.90691024629035, 264.93040508109783, 260.4716580044721, 260.15091461127304, 259.7344605052677, 258.24563919564264, 258.294123619139, 261.68880838252016, 260.6832845400784, 251.13676283904425, 249.5232973049575, 249.60093451010172, NaN, NaN, 24.0727244341814, 22.927237438012945, 22.812792251651622, 23.582489533614897, 26.37786644936893, 29.618045581211504, 32.15489866775855, 33.03293900739191, 33.249799203666676, 34.643597002668606, 35.59302550465388, 36.90852855086038, 39.77104622003405, 41.12808982149047, 42.998655897969584, 43.5458339315757, 44.01823714129272, 46.07106047162932, 46.35684916473435, 47.30577416833734, 49.76166461392097, 52.51316711756954, 55.26300195520225, 57.82692451079813, 60.394574695384044, 62.40776348619432, 63.51045478561535, 65.1601796669838, 70.2933030432763, 75.43075262885728, 78.35550912266494, 78.54040241137947, 98.53755356537876, 116.14489651216925, 122.1938781956997, 119.62963761050251, 115.77431454163995, 111.5536418779491, 107.15308972234497, 98.88884470465707, 96.98308554936816, 98.29802111807386, 99.6329130753362, 103.38331208751485, 110.87916411436464, 130.30564241282312, 149.0782031561584, 158.17956162181642, 161.13333213457778, 172.0333079119589, 176.2141800222872, 191.3673850766283, 215.22335522326003, 227.49963505497175, 236.01533911089697, 243.1338886888602, 245.44700329764288, 250.846582580548, 255.56915346064594, 263.12296479913834, 266.2548605492832, 263.09900017683304, 260.23467543920265, 259.2744369859988, 258.2219624856614, 258.1620986601019, 259.95976656886756, 262.76695111991495, 264.73013668996964, 258.24560405403986, 250.58080342842757, 249.79723311555622, NaN, NaN, 25.762190882655815, 25.831559043501297, 26.161642717841158, 26.30292638654613, 25.820415498386428, 24.967377384541606, 26.508767367090588, 29.120618804037232, 30.184429250256407, 31.797498366875327, 32.19684620564841, 33.88463924610451, 37.74504738312496, 38.21948933865047, 38.32614385392236, 38.91215118240912, 40.673726437258935, 44.12725709461457, 45.22366111344367, 45.73451537772872, 48.00896435697227, 50.20891280929631, 52.223568600069484, 54.976278462864435, 58.093449004436984, 61.210420763464846, 64.5061515021554, 72.21198488091675, 76.06705013022274, 69.09161508882573, 70.1812748688335, 74.21178017121606, 81.91303636333635, 91.99604047294125, 108.68841538706033, 105.21394643995254, 83.56142691179107, 76.39599721738522, 81.52876474647711, 87.94418361522578, 88.16518102262563, 92.56089527154451, 103.03685292213922, 117.72650527670116, 137.39036129620527, 147.8919274585491, 150.5442042378235, 155.9048299113575, 161.99368857827963, 168.88205284075948, 178.03997450284652, 188.821513146362, 196.65316421783325, 197.3615682006672, 217.7140037205315, 230.54570770418258, 236.54731264730304, 242.37210081337133, 247.00603187977038, 250.65561877483395, 254.7196410481793, 261.6869690589768, 265.03436773937375, 262.70588036686513, 261.2563551451896, 260.48803249644294, 261.7306400197147, 264.61495423269236, 266.73085038922665, 258.9351282767385, 249.96917794500695, 249.48139961917767, NaN, NaN, 35.30825020478774, 25.129951113653078, 23.688906658773146, 23.353516038622463, 24.233708560587804, 25.776446092523408, 27.758309961138913, 30.510688031126094, 31.28016791318423, 30.72218723767441, 31.59704809413307, 34.13002674374617, 37.98724279778109, 39.74835530636041, 39.08182085442814, 40.28303040334022, 39.950759186814466, 40.05314659466238, 42.36101709296879, 43.680855806603525, 44.88491095409516, 49.17764009154527, 58.53281194589245, 63.59388581796492, 66.45561787252392, 67.00629991785202, 77.25299324176761, 78.79232101881736, 81.10225126707408, 83.29877409506301, 82.30578423428918, 86.69815250795796, 86.69711801920509, 81.18627210488162, 70.39293028133764, 68.07012220460251, 71.03623374414869, 79.83692205316133, 84.90321408343763, 90.1886422408779, 97.92589259304084, 104.60584003957936, 121.03804889004289, 128.49517906021447, 133.41533893281073, 129.57718807440733, 130.65752585703552, 141.52257923413285, 156.24971753250495, 168.1796833204555, 177.85188709547526, 181.57374898457815, 186.13994752488034, 214.69122551569365, 230.7657015926468, 234.80215652710444, 242.82194606272907, 247.59111969033708, 251.29422167084564, 258.50230560345784, 264.86643896383566, 266.6481752197208, 261.98691515907666, 261.77109907486476, 264.34558207782686, 264.7403465570867, 266.9385840749869, 257.18217405298475, 249.89280205932562, 249.6305030010472, NaN, NaN, 27.26170989747274, 22.46520610118275, 23.051145591986288, 22.608992975694175, 23.563595641961847, 24.372930087830884, 24.88532601761918, 26.28117602060563, 27.60249446935944, 29.73236777294117, 30.75936920295108, 31.273596817459055, 34.50651020303616, 37.81578910224532, 37.29643365060632, 38.24347078207236, 37.57515589839194, 36.101778921784025, 36.53469677803245, 42.03877908438102, 50.378091907046674, 58.644514442596794, 59.97017250680862, 62.38680455692706, 61.606135232356074, 63.58022936367637, 65.89085907128326, 76.80022344404112, 80.98088366928522, 83.84036675777968, 85.93095970904803, 84.60339991514839, 81.85044254173106, 72.48149038438127, 65.31367461626475, 63.652052712432194, 67.39542195722407, 75.98127229503079, 76.96877855712314, 79.71548811047231, 88.33588148588916, 108.88229697515992, 108.37680478833659, 102.98724874410593, 97.34310985954926, 98.37812479515203, 103.78517399794927, 108.41358089530266, 114.58946235746845, 125.41114058943676, 134.19503001575112, 138.86585945406253, 154.91317083383578, 157.3716388788542, 162.18762420188781, 178.39709027221326, 209.332270177207, 233.0317480848918, 239.66680999189606, 248.38706686549102, 251.0445948109897, 255.16421875491952, 258.9727143943467, 267.3138989598365, 268.73042936734765, 267.79904365290196, 267.53764073077787, 269.69792541827314, 265.6263509555531, 261.0496341618981, 261.4152519456078, 252.5351262817969, 250.16005265005577, 250.21952440687133, 250.41756918571144, NaN, NaN, 23.88434330649226, 23.14482445536396, 24.321541915308156, 27.11500330012194, 27.33489574556495, 26.667104414630852, 27.39788726689347, 29.45586863519722, 31.439090405073426, 32.46788587304068, 32.979431540934264, 33.86088603617654, 37.6796763071438, 42.67939396358457, 45.105566121907145, 44.218134010676735, 46.04922067793976, 51.92320958576213, 53.389162740563606, 52.3550685883428, 57.786823016790734, 62.045434449675795, 68.50893824363644, 74.67619605811475, 80.55352861296099, 85.54715938336471, 87.45082105779704, 85.98047928691186, 72.90268522669643, 64.36145263275591, 63.769482789943986, 68.90168774136633, 69.18294205481712, 76.67181552603348, 92.67218876854312, 104.11817605449447, 96.64232227604214, 84.1673660951171, 79.16335058198722, 79.73596763342088, 81.8123145465582, 82.68760305555156, 92.385448891519, 107.9923164914636, 116.22187489069945, 119.44342506376331, 130.37082959875931, 141.60109334785352, 158.45886077012082, 160.6732937163886, 167.93925483829423, 190.6303072481097, 228.0703491796044, 240.72860419866944, 245.86461892797715, 247.7116158940876, 251.97418375224726, 257.229904481269, 260.9904867738818, 260.885315748859, 264.8057775764541, 269.0830615041803, 268.74087053168074, 268.7565802000839, 266.2704885531855, 258.83070336013213, 250.8836178546742, 250.37346437980062, 250.482188134422, NaN, NaN, 26.91560119118248, 24.922600459704135, 24.992473926522248, 24.841792072737388, 25.722161525785236, 27.34022359403961, 29.54745005118419, 31.23628505614469, 32.777707340919406, 33.80365038959245, 35.26994103176784, 36.29227772743999, 39.52511286817809, 41.72544065496074, 43.40743676445002, 43.69721693397337, 42.808757170501224, 43.83369771023844, 47.06163671209357, 52.2743863966181, 57.38004130757976, 58.91767449669858, 66.40380625692119, 74.00488086978427, 75.53900327725971, 76.63876853968644, 80.93161573001429, 79.05031014801108, 78.38516137695167, 72.76679802255008, 65.49092076155529, 62.618419412352274, 60.62725435613878, 63.7080949834932, 64.47662222544768, 67.3299635463707, 76.12911102211027, 88.7863452119762, 85.49444733382211, 79.20187708300948, 78.3434139501256, 82.74336788208531, 86.04807324234315, 81.64153203448647, 82.73767674374506, 89.13076940026527, 99.95741223608537, 111.21853834099889, 115.61561552821925, 119.36559230247028, 125.33683699491165, 132.91763112737988, 144.4785133279802, 154.31516911191295, 162.84315715470703, 178.4276511072714, 204.4911317377362, 223.45085300630498, 235.38511793726622, 241.98811400708192, 246.3704989839322, 253.4918276124097, 259.8390585518896, 267.10316950133887, 267.09659129126186, 265.4524510524574, 264.228255142906, 263.0642690571049, 260.44649697002797, 251.39618503960176, 250.23466442010962, 250.4034140219021, 250.4815077276214, NaN, NaN, 25.358737384365874, 24.322425104548515, 24.024396771886043, 23.946449720857693, 24.531633605060197, 25.7801701579695, 26.143493527799922, 26.652771247170246, 28.12142313187899, 30.02905256194886, 31.42179499571172, 33.40477086007299, 33.62495972716489, 34.43401972466389, 36.12278552022371, 36.855064291611654, 41.115451532578945, 45.96426496740814, 47.13685963821172, 51.69011269455098, 53.96583077649982, 56.05388787072498, 62.77001659844596, 73.79436882263947, 77.421562906021, 75.98503243024165, 75.10906683320577, 68.39103641154715, 63.53741532221001, 61.00515827621207, 60.1163799785359, 62.31709027306107, 60.7645166710204, 63.50780270765836, 68.68032396547498, 78.70591433411823, 81.45498169735504, 77.70459655250909, 76.04208848300443, 77.46168222567714, 80.6856721137854, 84.20786948360424, 82.01400266523117, 83.76575539748268, 83.99133167374309, 95.67355019942613, 104.04477765537978, 108.22859760455201, 115.94123791616003, 124.34413255609972, 128.13151077636056, 136.5620051909728, 149.22774945227636, 160.56719948554553, 168.22181084640627, 189.43577244283603, 217.07796085212445, 230.51900366017725, 238.6442847261904, 243.81672482189052, 247.59844726742253, 250.9363627062154, 255.56322048811498, 261.0311370458273, 262.7888841756611, 263.1376970590292, 263.6951721401736, 265.1467516650948, 266.12727065114046, 259.53311375630557, 251.26949066907696, 250.2749580161077, 250.45169003642195, 250.6229396826448, NaN, NaN, 24.57333480973295, 21.548979361961326, 20.734445154943487, 22.05399651465205, 22.199783333499354, 21.899397303398615, 23.071140672510683, 23.951780593802468, 25.346128431197336, 26.152421601263985, 27.619764287491307, 29.750011745090394, 29.821873919348196, 29.155119740274476, 30.47727888532723, 33.566864679159735, 37.97426746259373, 42.97081014766689, 46.862808309241856, 49.135146645989266, 50.634028082948525, 56.91019178065363, 59.22311493828009, 61.19786844401289, 70.99981119688033, 74.52427341105415, 67.80933982650546, 60.86299760459404, 57.992861172573754, 57.663771757706435, 58.98518993009537, 58.425819516424546, 63.378176269314174, 67.8860222201202, 72.3887234546122, 80.19948055408382, 83.82994754334838, 79.8639225441429, 76.7655582983192, 78.07641712867618, 81.12372534109157, 79.06873222857374, 81.11988924005558, 82.57704375503818, 94.02152654901978, 102.69728668300216, 117.40183390563632, 131.43389542356257, 134.86780142280725, 138.88207415642344, 148.0615649247149, 163.312352735002, 176.14452285233878, 182.0580967151739, 200.1362794617418, 211.81153451012977, 221.97225301976445, 236.89947703919785, 244.52882008584828, 248.3670226974487, 252.79900859104245, 256.15771341430155, 262.5633403494601, 261.79524199899106, 262.91152741898503, 260.8422486246824, 256.1134496458867, 250.8078255201605, 249.98928569365722, 250.24311585159066, 250.49104608029648, 250.6124541302421, NaN, NaN, 25.71861079808457, 25.569194720506815, 26.007908269036367, 24.08953510835175, 22.83198634354273, 22.46131223334869, 25.625842358317332, 27.906339821455038, 28.490439901630655, 30.326313492479148, 33.635540845453676, 35.98412273144104, 36.34833466259014, 35.460782174689356, 39.13225873732316, 45.010364751012055, 49.78562334215276, 50.88864883371632, 53.67217143313281, 62.261445403468805, 65.5352340777875, 69.279805984127, 72.24580340792403, 73.6696908522273, 70.91442592698978, 68.04442385909418, 62.6378474584535, 59.329137681787266, 57.996127241851305, 59.52348377546369, 59.40145039750742, 58.62274715511832, 60.92670798337209, 66.20228125814494, 72.02872910876872, 83.58276967854606, 83.26564194028859, 78.96223492425163, 79.51006165970288, 76.96861422038278, 78.71798233142938, 81.06542694809264, 95.33221554604329, 113.71616902813012, 129.30985543627153, 133.78337099041332, 133.92966449343214, 138.52942645928727, 146.39245472232676, 158.13713072688725, 170.99754282403242, 188.98626621601647, 203.65936476361205, 214.52454289971766, 221.8039699647954, 235.77646736362783, 250.49089795482843, 256.6904580258962, 263.82681908564814, 267.3008004783897, 265.21935459551014, 265.1214492029418, 260.69563716998124, 257.06454690091556, 251.20374492699045, 250.30280024640234, 250.34642288618667, 250.59592500495842, 250.70356520767805, NaN, NaN, 27.533460915202905, 26.941568597380883, 27.30827140181719, 26.718361490899017, 26.123774494961644, 27.519751631209406, 29.35568186491634, 31.4871943930944, 33.98897329572372, 35.8247983184948, 34.05227670252315, 33.52668005845386, 38.743464125385806, 43.298335504482374, 45.64781636958496, 46.08167297553537, 45.712007653755535, 48.721967355360654, 52.9061922725602, 55.91531943570197, 58.739669041795445, 67.21499380590518, 75.69361232664698, 78.21960509906845, 81.30472661075268, 76.90180719097796, 65.98024399864923, 62.00910514676556, 59.46603912820948, 58.135041757836, 62.098936867329655, 66.83469804078257, 67.70445543993031, 67.80228962738174, 71.42124698011125, 79.11748924965976, 81.30233646849123, 93.95433278644181, 104.5135396733859, 93.39475855394537, 83.768571647576, 83.16765548860562, 85.65987124998365, 96.98177077493041, 108.30724903481897, 118.61204102677367, 129.81771973184956, 135.0211664798789, 140.06730669663222, 148.05833488987003, 156.52467046273688, 163.12959685295957, 174.3024608019436, 190.8539597859471, 209.3768670718783, 220.31822921717563, 231.52530764653199, 246.75766528139567, 257.7852843374975, 263.01602965433807, 265.1549362997359, 268.3055510381424, 263.3666842125615, 261.30645724028744, 260.3110368599979, 255.04408066427197, 251.2950092974691, 251.24161466569484, 251.33958416848725, 251.52927584690391, NaN, NaN, 28.488830223310902, 27.78526577421582, 27.782620447681772, 26.748322918019195, 25.381585404236628, 25.56230538431408, 26.072995115279536, 26.951808602548446, 28.56884249552694, 30.84722296374806, 32.4585073991326, 34.47681132213093, 36.606138199130605, 39.13822244535237, 42.36949681431979, 45.41182999269186, 45.33373458025762, 44.15324122721631, 44.80501286204341, 46.413662708806555, 48.83394662696401, 54.118402448351496, 60.28770789047094, 63.25906460224695, 72.73354335482395, 79.34227084057396, 80.66137047907233, 76.8144942008284, 66.78626251537858, 59.0627290935619, 60.158550327675044, 63.45971820568462, 64.33582799399518, 67.40944432767861, 77.31722774569504, 83.47460407250298, 93.69949788936563, 103.04355670550517, 108.76853781057535, 109.63068428466886, 109.84676673485467, 109.48591931030205, 109.86239156763558, 116.84080004219044, 135.39978697571175, 139.4578757966158, 144.08789821586856, 156.4792504347996, 161.65010970116543, 165.9392878441992, 172.14055137514336, 176.7569200847676, 183.5210967567008, 195.68126387302073, 211.98912096990634, 225.53798834825966, 235.72280535194068, 248.877876103186, 256.24372878899413, 264.5544619114352, 266.8770267811223, 268.0184391378469, 264.9437278918893, 261.7374171988447, 259.6734338730505, 253.98706765973677, 252.39132035552288, 252.35935502897917, 252.59247315145006, 252.76135701424008, NaN, NaN, 24.692477012286624, 24.17443519955296, 24.39305697646648, 24.535155303123055, 25.5614001426415, 27.325478485023616, 29.01465602872216, 30.40798283923788, 31.72908085819345, 32.755357532091764, 34.74143754944587, 35.1779964844333, 38.0425324220817, 41.345416141659676, 42.29438286080566, 43.09840643625523, 40.15106929772378, 41.09447493906094, 46.23128260333676, 47.69651859581552, 53.53177767976997, 57.20421261867309, 62.19438905388529, 69.53247494731717, 72.3130518425961, 75.09261492923609, 75.5283049703107, 70.38172613376813, 62.7463518429553, 58.3335825342254, 57.74038418754818, 60.6727780190682, 60.510191351014974, 59.76828078016057, 61.67015827604925, 64.3015096281405, 68.26331777673876, 72.95612942019902, 85.86632981026268, 101.70739225204416, 110.19566378808854, 110.5095330440081, 112.71094029890992, 117.2277147877869, 126.02208124256751, 135.3052195394126, 145.9051546463941, 148.66850690965498, 154.45425499588347, 160.5925177157525, 167.25059627570118, 174.5334413869418, 182.93615162102142, 192.25149182253972, 199.40534877537218, 212.07374624673346, 223.03595056404353, 232.49936554983367, 245.02772292123183, 258.1722750579602, 261.4587000068985, 266.37064388771654, 267.64397257806803, 265.6363556059804, 262.6564719603934, 255.9248696233205, 253.2033540748458, 253.3737034084784, 253.62003879271532, 253.86524428614428, NaN, NaN, 27.310643300716613, 27.162052680602137, 27.52659839730174, 28.40750095896439, 29.434263079283284, 30.460262453415233, 31.70969100103532, 32.883870177329555, 33.83823452588859, 33.688920416745574, 31.329637222752485, 31.615793441267193, 33.45305762833466, 34.10656238836679, 37.04298897072282, 42.554181197706896, 44.463485376207295, 45.48637983128707, 44.379579544907315, 46.87366769790355, 51.57116920054635, 53.91961072111926, 57.00021647604801, 62.42956030755495, 68.66789498023695, 67.63680883372749, 72.55324788113366, 74.8276662718009, 72.02899927344613, 67.69643098413768, 62.327425521942274, 58.06043437473299, 57.02064421410005, 57.30428855797124, 57.51908051484363, 58.980910000547176, 63.968693102719705, 65.49911506573805, 65.92905146035149, 68.93317303237743, 74.60668497119346, 77.16388961323283, 79.71919500949751, 98.42168385573554, 110.33811834828064, 112.72965537913328, 113.452307480802, 120.42400150497322, 125.37248527559582, 136.79253726861913, 146.5627172366468, 152.28473652829533, 158.62802338265294, 165.89742074234695, 174.1048384841217, 182.46853305850627, 185.8645435040806, 189.29267000389845, 189.44864785650577, 194.6655062929321, 208.32056239376092, 223.09149250323225, 235.2556803711234, 246.2229342264312, 257.87847824887336, 262.4350730048002, 266.5213978811549, 268.4181143488071, 267.00507659366735, 264.4155672513499, 258.11543841568977, 253.69259266518372, 253.06188543084144, 253.45467551431975, 253.83615139910864, NaN, NaN, 28.350335901182316, 27.831690477242873, 27.901907299881284, 28.263092836948296, 27.962263718710656, 27.36633488913661, 28.100200630963684, 29.051999033042353, 29.488470819047535, 33.53173508524333, 37.13378683294288, 38.74739623098189, 36.97873745137939, 36.162675637783536, 42.33513990567928, 44.31469903148261, 45.853365410531346, 47.24345098534224, 49.6625453518759, 53.844647056249656, 55.088087114310156, 56.94749279950282, 59.80492535833794, 66.1913133354376, 75.22238811249677, 79.8406074254562, 81.6988260994737, 83.01478593292163, 76.40909363922772, 66.49409770470342, 61.97867376670844, 60.761008220157144, 62.8430892413488, 66.02253665332488, 66.56001233657325, 67.98028702260723, 73.14297144207956, 84.02296518214233, 91.16717123655526, 96.01295003450264, 105.79413989315886, 114.16982585140039, 115.6432017934386, 119.02297751100633, 126.23430738662752, 144.04418311005833, 151.7276548039059, 157.39317275765944, 162.86422645564394, 167.7812426644674, 174.9338909124586, 184.32030710992268, 191.95051211535574, 196.2922402677783, 199.66266841408083, 213.0947510998565, 223.62120576929394, 234.4414793513058, 245.65397135466537, 252.86057952812553, 252.58020110326999, 263.8270302118544, 268.48005931353964, 263.1270223986873, 254.64837805790415, 253.31222737899728, 253.0659953957634, 253.24975637432743, 253.42052926497357, 253.57970290634813, 253.65152366421117, NaN, NaN, 22.84893112811097, 22.256798261682732, 21.88466682950433, 22.100441390580677, 22.831995852368554, 24.594516843905662, 26.282723054091978, 27.16393854278461, 28.779141471968757, 31.05861272542491, 31.640470443265208, 34.42974992917273, 39.94070738216074, 41.698315348956555, 42.64689640324531, 40.737143995615234, 42.496287914925446, 48.15085464972868, 51.08364990627904, 53.21162993246123, 54.0873618762045, 53.41771471610621, 58.2637154694412, 65.85663412725451, 69.58945568983526, 74.20876513293915, 79.26432485046512, 83.22572083439773, 79.48531443107714, 70.0116708667731, 64.83014211637904, 60.19749074484268, 59.521769027091665, 61.381316223207044, 64.44969971715831, 66.64467359177014, 67.18797162963791, 70.81169051406799, 82.03048080500434, 89.29195555836904, 103.47104643305262, 111.88567557569081, 117.3752607780055, 117.55790779247774, 124.3875373192841, 136.02818178741387, 149.13306035960966, 158.00909690636672, 165.80794291056202, 175.50607004320725, 184.05900943191878, 191.34271730816235, 190.5345817428972, 188.21791187355353, 209.6935198023795, 224.5336971137796, 233.2710848392783, 240.57524555446423, 245.47547644742357, 250.67125559775408, 255.50993440680043, 261.48283571882314, 267.0057828646319, 258.4322565513611, 254.76956307718822, 254.41812288336902, 254.5151202932451, 254.536435153755, 254.511239004087, NaN, NaN, 24.357282523823653, 22.992904794951418, 22.179946007433646, 21.917885029694173, 22.281954084976867, 22.82871716584385, 24.223186805490993, 26.208231150659483, 28.485881017730012, 29.031771923633563, 29.653721503732065, 31.635272643472188, 33.47175340825267, 33.317441066730616, 36.87844237282966, 38.64050376934245, 40.58427222264477, 41.351695193969135, 41.12826865791851, 42.44357261855544, 44.20251663454645, 48.381355812495876, 53.99972257230087, 55.645881441709655, 59.16387159821227, 62.79520294663963, 66.42119942320292, 76.000516661827, 81.7245942853368, 79.18785616005643, 68.94439599486778, 59.9038439942953, 57.577661710643355, 56.908257299807616, 57.89243189524782, 59.53867220935293, 63.27193041153282, 65.68197364671417, 67.4349399986525, 68.96972916347036, 79.78638650630602, 95.33680134662491, 103.41414789175583, 114.43153666743477, 119.14026631617698, 122.80919581865002, 129.57633743531295, 136.79761049927586, 142.81858125692284, 150.66904123614842, 159.43072335111435, 169.11842141872324, 182.67966386464053, 189.64827811288887, 196.40938744458452, 196.51692074309713, 202.04244899338642, 218.90920689588586, 228.73314346113037, 235.43290685350743, 241.56099050466935, 246.58713105983563, 254.84488240894356, 258.07332768878535, 258.05730956148074, 263.3977701523268, 257.56146534840644, 256.2969446244714, 256.3159700592827, 256.4849955877642, 256.51103601603046, 256.39682088763027, NaN, NaN, 24.511126677968452, 23.881433106762948, 23.806607643648697, 24.318624024284304, 24.534949637853657, 24.49273071340065, 25.555760478673083, 28.278699070226494, 30.15182698999554, 31.434704515483517, 32.09117186601039, 32.04902726615771, 31.640861942829353, 31.964436401379913, 32.54737608624166, 34.56435498799286, 39.00830737396652, 40.06942360293939, 39.547267588952465, 40.79098861895026, 43.87554103199753, 48.57286043781515, 52.68099323327846, 53.33969668173592, 59.504220851609105, 65.44450023189748, 73.29786897732572, 78.73246511461205, 74.24912730897633, 71.37510878830518, 67.3351880131362, 59.33061716947657, 59.32627206107298, 60.49606717374317, 62.02919000622232, 64.88353620563572, 67.22584864281386, 69.05331111140221, 71.53884357130401, 77.25035013894929, 87.3659672264713, 97.26252768456929, 104.31098912928061, 114.90646037057518, 123.08272285298591, 129.59210400556432, 134.66629129486617, 139.72753292742186, 150.1677101941871, 159.17100139934547, 164.63836295711403, 176.15973825606488, 183.61199580515935, 189.52285635950957, 196.47838046325458, 204.55803203181995, 207.46829982784703, 209.345277416351, 219.5654654565998, 228.62684669969764, 234.9268414640028, 239.88875065743596, 243.54727757067397, 249.91696811549227, 259.49350480389944, 260.8173476002164, 262.95026699042046, 259.37727564248075, 257.1365548927822, 256.9809575292073, 257.1568650121858, 257.20522340887914, 257.28915785165674, NaN, NaN, 24.99274795906107, 24.473008361135932, 23.254630397023394, 22.698137337749994, 22.87937974629056, 22.616320855422693, 22.9799585979357, 23.600291522547437, 24.55147679419287, 27.858872561500675, 31.832933039367923, 34.331881937684486, 34.17893127859248, 33.88193841749157, 34.39258195552155, 35.123910918274476, 35.74245688318862, 39.52099730438627, 42.01831440517978, 46.41788641527372, 47.04221120621343, 49.682495978690746, 52.87379806926168, 56.61297788068344, 58.58891182996236, 60.233001453294236, 69.03721657610498, 77.5102357954179, 80.2524626802618, 80.79210622254666, 77.70440273698355, 75.3812179328171, 64.37921090238036, 68.44205437675708, 71.52094835466876, 65.02042107064521, 63.259553440258465, 64.90954409859226, 69.09021664173615, 74.58609705960447, 86.91702058314222, 95.50051045909676, 106.62480382474723, 118.7377857259313, 124.45958471290207, 129.3141367246454, 134.51225381870802, 141.59337824476748, 150.78651833634248, 159.67522826261677, 167.15105443435692, 175.41249007482077, 183.78093854775628, 189.90607895201424, 198.7893127357174, 208.19196182022668, 211.48404824271913, 218.9794686011327, 226.17433991065266, 233.03115242771779, 239.9218854648884, 245.62900510844813, 247.76889495660697, 249.0573198609007, 259.2757274767783, 260.96416268279967, 258.8632609982989, 258.1774080487945, 258.14244860431734, 258.10257883946923, 258.143049849519, 258.20581572124075, NaN, NaN, 22.921249991581494, 22.698089878114573, 22.91862490564805, 21.84849228863081, 21.84380843010252, 22.206582819266394, 22.642180757637604, 22.892857683889133, 23.475442735087377, 25.34445031643616, 29.23865600973476, 31.9205435956686, 32.62071116555306, 33.385368471497294, 34.85298587666026, 38.23295132344944, 41.537353408001316, 44.43397820866821, 46.59631461830907, 47.21845398337275, 48.57133390362745, 49.557436842766975, 50.87737011984542, 53.07482805719801, 56.15332170242138, 59.01456564701947, 65.72213303216483, 71.88392800482322, 76.72312488865867, 79.02478450239843, 87.93695755268234, 87.27811425952399, 77.69602321550428, 70.08567606833874, 66.33733418702583, 67.43846951027454, 70.40634217377598, 74.69094609663195, 80.52712766354954, 91.09843826797781, 101.8324998863108, 106.57272178884277, 120.31727096905543, 133.7785095854695, 145.6218747285753, 156.08664499094564, 164.09899943001463, 169.63743568289522, 174.64119147326252, 181.03751619780675, 189.51863685152583, 198.05729855560725, 208.10706235974985, 212.69854460453647, 215.73305466099706, 224.53342132332955, 234.26886186348688, 240.78981483547955, 243.70271425917852, 245.36516161641777, 247.2164834705218, 248.40572837406415, 257.1412575985613, 258.81491554318296, 258.55839968261864, 258.5980444561154, 258.83142488394384, 258.86107774888416, 258.88014499154826, NaN, NaN, 23.47984732846323, 22.480282673190104, 22.549989838052444, 24.01713339056333, 25.560135626969046, 26.364738394662695, 26.801433657757215, 27.753160978847827, 28.703168285506624, 29.2507254441888, 29.465311626354076, 30.15673068462509, 31.25312193707472, 34.48077104527635, 36.35037964698875, 34.87490977658758, 35.49487704240066, 36.81038271151353, 39.4135848399054, 42.091911680112844, 44.3641895374533, 47.222735779324374, 49.057634125519044, 51.40087609875579, 54.11237997639965, 54.913198801963205, 56.006765839879264, 58.20457412335113, 61.93858772473933, 67.94904940391393, 76.38630327821812, 77.85824293658355, 77.26728856392272, 79.98022460234819, 87.16976658218586, 83.49706629264786, 83.56682522024391, 76.58646778083073, 78.56220724173691, 81.63162943617674, 84.27793270997337, 92.16407850075726, 98.96195631988783, 107.04334377419035, 126.85881454301501, 142.48559383651056, 152.99794244775725, 159.30746878500827, 165.9983463798146, 173.6222561257817, 182.0189997060376, 192.66081505388223, 201.60698342575432, 211.1855123317728, 220.20078700078264, 230.31342545511063, 237.8211748577448, 242.63277501471384, 245.50580270172424, 246.30477778776708, 250.1839449315605, 259.7083630837701, 259.31808319921834, 259.3673711214051, 259.3199940487923, 259.35084342073134, 259.4483158412292, 259.47500253005296, 259.5153539638373, NaN, NaN, 23.76866838295542, 23.39901356583037, 23.101518917319016, 23.170932990069222, 23.38870252722035, 24.121347894064897, 24.853309865878654, 26.689849419539176, 29.191363882659655, 31.100802299740575, 30.950025013005746, 30.945503806764055, 32.33827730299733, 33.80218977824396, 34.16467769617941, 35.631901936246685, 36.949654511869205, 39.4404324001899, 45.609642558289, 49.86565305865479, 48.06369256360534, 50.85173273025044, 53.339056354086956, 56.05131615240725, 60.81937337215442, 63.08857216419796, 64.32893365201528, 65.49227167862013, 65.77656324705265, 65.69149021975463, 68.10797545867008, 73.31232005002691, 75.43878384132634, 73.67096379008329, 75.42851358624058, 78.72076709181954, 81.43050337316427, 85.01083053217475, 88.3837653517951, 94.03652593622284, 107.92596261184785, 117.41721688972538, 114.34630228727545, 105.12263656358913, 100.49960948031337, 109.76793304680977, 107.2207358818388, 105.44855354039125, 122.18243510650181, 153.62729466466013, 162.92292179133557, 168.63403081913472, 175.6865622422391, 184.85203542931302, 194.77120997079948, 203.15418617081673, 209.6194722190849, 217.62006135670444, 221.93764325015604, 227.45285227844136, 230.38822212687643, 235.27735703666082, 239.81468253952002, 243.4733829751724, 250.0370646406156, 254.06922007907602, 265.8256673143143, 263.17625909670556, 260.9403164822057, 260.26986462083454, 260.018804974935, 259.97307806074815, 260.1642315282826, 260.36162256443015, NaN, NaN, 23.324871606394634, 23.912974285262262, 24.057492132839222, 24.56921065207739, 26.258326585943994, 26.47569101096354, 26.544157315602504, 27.94059361936477, 30.07041510677603, 31.75967222889296, 32.49271604679661, 33.8874190727625, 34.98477297520485, 36.964052548811566, 36.95840688707587, 39.74751773191669, 44.66721294243368, 46.495402376366094, 48.174283004878525, 50.815324991622035, 51.990298631394815, 52.135385756804155, 54.257300966127126, 57.33906996150267, 61.891397664883606, 66.14872593217251, 68.19869530465988, 68.62980933847311, 71.92752122161923, 76.11054189582994, 78.6682263330446, 79.61263324141494, 73.36994717942741, 73.06521391502184, 74.23157993950247, 78.03617867611821, 84.11904950760947, 88.08501870063628, 86.91430292866308, 84.19560925411855, 90.0602159597067, 94.90264890291819, 99.74748317938398, 113.83900221498135, 118.68803134549951, 120.44308477264816, 116.49775368564748, 112.55166359112452, 135.9126851477862, 146.96134239641748, 141.5353075517272, 155.01190854618605, 172.53826534479182, 181.00364661265104, 189.04204213056008, 196.9135039843079, 210.21406207652626, 220.45232434401635, 223.97818515891572, 227.51410494020706, 233.4514231494166, 238.99929179011085, 244.15180762133704, 247.49333632084418, 250.5594512702776, 251.47749375858163, 259.63516741903334, 261.3289905939385, 261.1898117912764, 261.44237081344124, 261.5345655722312, 261.48829742703464, NaN, NaN, 22.372350948037045, 22.442969757441546, 22.365942078394212, 23.170493410809126, 23.756057798729394, 25.29836936331491, 27.13265407998068, 28.74555432688957, 29.180669459226667, 29.836132680071167, 31.081491259256598, 33.06381499845015, 34.7536656950154, 35.704337508779254, 36.72885358994344, 39.36959763256427, 43.111891700175484, 49.425393028387816, 51.99267839726491, 53.604263126656235, 55.29146135888941, 55.28100133269244, 59.13112883038762, 63.20129697329753, 66.60933520516527, 69.35692440623644, 68.80109431582355, 72.31035164145524, 72.96866592936499, 74.0623510801101, 72.95801238610316, 71.85462609360853, 78.6797319999622, 80.87751761957657, 91.42807727287378, 84.05069794077943, 85.3713389906603, 88.66531714310062, 92.50501877516751, 95.25829719807423, 99.59446904702226, 105.97666094229466, 112.35740200876295, 118.752722052431, 124.2711266928087, 116.60860933597695, 108.68006490910157, 111.55879771164915, 125.03221554855429, 146.21927203700233, 170.75299627260856, 181.43340053273604, 172.75117134342278, 185.2165189355785, 202.2177353042708, 216.62608734774298, 224.48255776414743, 229.58557934951665, 236.463288564154, 242.40409937008437, 246.15625550602235, 251.59561159597624, 259.60669590106403, 261.1188553575935, 261.33586569139436, 261.2324665768477, 261.4711801668349, 261.55931128266656, 261.65217183845203, 261.6311088541674, NaN, NaN, 19.42010680807298, 18.5678556575674, 18.601538372672593, 19.222900413231677, 20.248870378643286, 21.864308811434654, 23.29444729142733, 26.196070783360568, 27.8118896747558, 28.689309376801763, 29.270870634186902, 30.70212611588613, 32.20567837807113, 33.11905995287793, 35.20839306321069, 38.39974835404556, 41.296739300507305, 44.528065424178806, 47.24562474619134, 49.15249657914523, 53.51661233485068, 57.18039846903776, 61.21573839520799, 60.19410613789618, 60.18908880878852, 65.8379037636802, 74.20289121049385, 78.52633059806266, 80.64726319234953, 77.2752743146038, 77.70938849488087, 81.2210231897946, 84.51490895435772, 88.02066317339971, 91.60472147009993, 96.07814445171353, 97.02553494371269, 98.77477898492822, 97.30858110234033, 98.68774324979645, 95.26909537008594, 99.21527931923717, 100.97741323357889, 102.97025464623142, 106.93988782775635, 112.46278639037291, 118.64811778250912, 107.90374806180878, 105.5064574502367, 116.78234999145165, 136.44275910455178, 163.3977927940024, 182.75762318755687, 192.24150287342277, 201.12581641645346, 210.89947200445803, 217.75244568342123, 225.0970582200656, 229.1955063577124, 236.4241313274281, 243.0354829477806, 247.39056542439002, 248.82047221759098, 251.03241797470912, 258.2343775786146, 261.42309150807773, 261.9264470513766, 261.79536151250886, 261.8654058000437, 262.02437449640144, 262.1179119460688, 262.0011946476252, NaN, NaN, 18.96964206373178, 20.36598750302258, 20.953471806094118, 21.9060652036868, 22.48976156830404, 24.215425308824017, 26.23634782787562, 26.599209635160914, 28.948752076098234, 30.819125813012995, 31.95424690563738, 33.052272464017676, 34.84973650241402, 37.45669453821927, 40.02523076178507, 42.704617716214365, 44.4993652365535, 47.54561082853257, 50.80910305190776, 53.44969572915166, 57.705779147208524, 60.45083668065991, 62.42818710736117, 66.72100233493983, 70.57546594092112, 73.21429753784955, 76.39662689248149, 78.91655156628404, 80.8943508085937, 81.66337511850307, 86.28143121310246, 88.14595317108642, 90.88860028310145, 91.44756874757408, 87.04055583285165, 92.42329891287143, 104.74602429198565, 111.34015649266702, 113.31778782230171, 113.33646768286367, 110.47768542447392, 113.31725697101783, 113.31109463216748, 105.59571276589324, 101.48620262187542, 98.92523306116979, 98.41236648114078, 104.61089061503779, 114.63611083347242, 123.89757015424843, 136.2588178989134, 155.9085750646204, 185.9358077876531, 201.78305224866975, 209.140644969841, 211.49770159720808, 215.35004865799533, 225.1365709505195, 234.31417981481493, 244.65744227768803, 248.61085559231338, 250.5588870037158, 255.30053995319963, 261.24840647472155, 262.01790745524306, 262.2651298631818, 262.4312894909976, 262.53435724294485, 262.56230070717584, 262.59674997072614, 262.64015436250327, NaN, NaN, 23.81138130630996, 23.291207819896744, 23.14074475188703, 22.766396510394287, 24.270895071232893, 25.48019923489026, 27.57189546998048, 28.26632587947183, 29.361688070573862, 31.08616370277941, 32.736825749322534, 33.465717528756365, 33.973321126313145, 36.172805788583844, 36.53783563664439, 38.003728427098125, 41.27196879839653, 43.213274688369886, 44.30864319805486, 45.32819986175084, 47.082753758134814, 48.83850073487553, 51.03129708977334, 54.11009616554679, 58.94962887650958, 62.24885928369741, 64.96455088656815, 69.14197799500147, 73.0959720507877, 78.15691993714309, 82.4770485250541, 85.47419380466897, 88.69681526354366, 90.98425838621374, 90.47324380794682, 92.66813907601528, 89.88638647807718, 90.54333026486962, 97.79429473438242, 104.02490883405119, 110.57166033498454, 115.36093982042227, 116.63504645862872, 114.81921700115825, 115.7597718486121, 115.21719010251608, 113.18776831990274, 113.01262035274564, 111.936073399754, 115.79318609085362, 127.39596817306987, 146.2190942681904, 159.33046901250208, 169.2884535156347, 183.39325484334717, 189.32760870821235, 207.1113001497939, 221.5226389513469, 230.90765747782805, 226.98273366963744, 230.61137440876632, 237.67152185526362, 245.60396593332868, 249.75851915289232, 256.4204146466065, 261.1440149451803, 261.6899556755165, 261.9373002319149, 262.0324480428308, 262.19217755124464, 262.21481478580324, NaN, NaN, 22.663871913186778, 22.144327975277683, 22.766452290562505, 23.499034136235895, 23.82661458176726, 24.630507800579778, 27.237516513894107, 29.700660724749053, 31.79281222697033, 33.10812173905932, 33.540113907129935, 34.30691241770752, 34.74308367046328, 35.69383870197674, 37.82702415584614, 37.82452475638437, 38.58981835418334, 40.86400323096592, 43.13845775955399, 43.20254755111583, 46.68800980440626, 50.1025112123604, 55.16257797797603, 57.14921682379112, 61.99325575885822, 64.62646497928219, 69.13105967763971, 75.18671747820974, 79.46979299888126, 79.24490095624722, 80.22695478372822, 80.66916220829089, 76.80875946683983, 76.24710536321525, 79.8605222858616, 79.86227501507362, 77.9817336199046, 82.15636424575956, 87.87946049785221, 99.20573579629647, 110.98312334943049, 118.91863102621787, 126.57713963077519, 127.92086105784097, 132.5160758579722, 138.2688836277309, 128.030682698218, 128.36703737339496, 143.40705969398573, 157.91456422978902, 170.50093760064553, 182.6947060509331, 196.2349079469951, 206.68093090892023, 222.98567232477268, 234.59309550424416, 240.495118902772, 247.15341865631967, 250.54872589186627, 254.1175007636143, 256.9059104292213, 256.1789892031892, 250.93307580188718, 256.9085628530457, 260.43584771442363, 261.28026328592733, 261.5931243741324, 261.6923516647656, 261.7220287301288, 261.91588745998433, NaN, NaN, 22.85316816738735, 21.779771056530087, 21.738142453817606, 22.32348098183599, 23.16560371460435, 24.48895461226784, 25.11004708375343, 26.615661409383485, 29.37222785302064, 31.943984185287487, 33.66779459501771, 34.84079845147203, 36.27119678707827, 36.99995729085926, 37.28531391272598, 36.98364095242974, 37.38184058753774, 39.03158268723344, 40.71364255766217, 42.399947148561154, 44.45525154025408, 45.18426957804029, 44.73771458352533, 47.95944876106829, 52.357079360068276, 54.186020323618585, 58.21957640430079, 59.91096239413448, 57.63166837034614, 60.042574290948366, 67.44437443930146, 73.15862917017365, 77.26631634130992, 79.24516704416628, 82.61851652690346, 87.60541960759464, 92.22577395288172, 96.62276188305654, 99.10911413648601, 101.9648600223498, 105.45254533375181, 108.8318280625839, 113.53591430539583, 117.64480703163221, 122.2015360968778, 124.71463966781648, 129.2877253854568, 137.2383672944192, 147.73128020281442, 154.0732993941576, 163.26853177843313, 174.85863809863815, 178.62800403187308, 181.98250031856102, 193.02749001250896, 210.44027573942193, 226.92820583592803, 235.2972381825936, 242.39001565711882, 248.01041342163714, 249.4916122102305, 252.99827830363282, 256.9571921907511, 261.3734880174168, 263.7513614006316, 264.9740997076113, 259.2708669213663, 259.1033364009283, 259.6447383102464, 259.88520471213917, 260.1975362121073, 260.44987688226695, NaN, NaN, 23.178818114345372, 22.77121107399562, 22.657121573173406, 22.323613178366976, 22.502104507662988, 23.712954976690174, 24.480197636770807, 25.543013399157044, 26.126669876052073, 27.631733215658983, 29.868119432622866, 33.06132622516403, 35.1562907737284, 36.108530823560315, 36.104755391605764, 37.27509291500526, 38.666710524923424, 38.21989117525577, 39.094972427584025, 43.167304263257726, 46.948552922496475, 49.00067826923868, 52.37232282807188, 56.11783952277293, 56.62801076846244, 58.60498202850909, 63.88497533808957, 70.19283867682589, 76.05240030035048, 80.66967257305136, 81.8290131258309, 85.48701224821711, 88.63023107156941, 91.03850287457219, 94.77223940280534, 97.77059313444978, 100.70811704960578, 103.5682240289593, 108.46750316754438, 115.72418134535259, 119.2863230920659, 122.42296361273682, 128.30662506780277, 134.374418657026, 136.78210335656777, 139.55985731194122, 148.82366451383348, 160.6652161067353, 164.0160791204732, 163.75037603850367, 169.70715071526388, 190.10514556318734, 203.02378828698963, 215.42027717794238, 231.08460417779685, 241.96919423312534, 250.690472688682, 253.6579011725862, 255.2684979682492, 256.2268302117024, 260.04482012620394, 265.0819776271921, 267.01743300416666, 260.5034614867368, 259.6089021968452, 260.449439195421, 260.9238385695786, 261.118955137815, NaN, NaN, 25.57685458520776, 22.070585558191425, 21.99493823928299, 22.61753119700935, 23.49844652953489, 24.930073942869264, 27.540608916692186, 28.567098621028443, 29.51923861964022, 29.549995262264478, 30.24181943561151, 32.924998936340906, 35.45908778480414, 36.481849531625244, 37.10311209346669, 37.31785540061959, 37.091670048012794, 37.85686496521483, 41.41672873926172, 44.24193555333553, 46.920273127329644, 48.384638891927004, 48.30615835456279, 48.222823059336044, 52.98873712683453, 61.719594161853315, 64.87408087425408, 68.8290717019554, 75.56758545769152, 78.33834700863427, 75.83884136176097, 82.93703931494466, 89.75063470079287, 92.89187296218962, 94.79546160728175, 97.28563233588716, 101.69188573639207, 102.94238196176971, 110.49583667383567, 112.55331742689319, 113.03774164114506, 115.23282524072513, 119.78224852822953, 128.30889149405263, 128.76165601610379, 132.03738663386912, 142.65152362394846, 153.7417730872344, 165.7540679414178, 176.58804548621615, 181.57331539107872, 178.51423969647107, 183.41263327201904, 198.2107396391476, 214.65599588527633, 224.09671830712932, 234.2416712683627, 247.1541155761633, 250.6881632881621, 253.23358122860284, 256.9046289333041, 258.3796120361879, 262.1163344914299, 265.5708565040498, 260.60461574197626, 259.98101783516563, 261.0461113749574, 261.8922006203034, 262.4437858008914, 262.41943475633053, 261.96584382346725, 261.54981415776376, NaN, NaN, 21.633954466596396, 20.45185652970635, 21.295512777565715, 22.508084317001252, 24.34472893715939, 26.184037528868608, 26.917859453627774, 27.76174272582257, 30.63103924580863, 32.13815073541941, 34.045467436465884, 36.17041545635715, 37.74383813786053, 39.541497668359604, 41.33458280482294, 43.16528906402056, 43.892949641269574, 43.00279626673263, 44.60840021403251, 46.43746640118443, 45.87993205303343, 51.16111129499943, 53.468052400949304, 52.57657664295905, 54.550048643919745, 54.21037808945532, 56.839902534443624, 65.08645981576636, 74.43094611172454, 76.95926763277544, 73.32661522456091, 80.57288917386894, 81.88435692523971, 81.99089967902734, 76.926690502253, 81.42220599048738, 94.05361189964404, 102.85289346098924, 105.82731526673969, 110.33119930444661, 120.3014713899737, 123.96034298558925, 124.62864474301873, 126.07684615668015, 129.0665246154337, 138.84431944681032, 147.57437428515374, 156.91388803732028, 168.72295425269618, 175.87361239071214, 188.8318743948672, 202.41896914015845, 211.06855613000323, 216.6348145108492, 226.07573504317432, 234.3697796877085, 242.43872433368102, 251.5583786193434, 256.60051181462046, 259.475324609794, 262.46385759429626, 266.22326167017235, 261.55027139276046, 260.37521384313845, 260.98913867237724, 261.61222668785723, 261.8200923993415, 261.18550258574123, 261.30898097941196, NaN, NaN, 24.36268434652913, 23.289345553634867, 23.285355670041604, 24.055384628318265, 25.745178812830083, 26.88318628095569, 27.356130417731745, 28.493984193176406, 30.551424327373407, 32.312648774014995, 33.99910666643657, 35.42728988998625, 36.30368454082726, 37.62127869609305, 39.41664796640294, 42.27998755906704, 43.30393286577832, 42.856808616751266, 42.95856604368988, 45.23314884617674, 49.27336939065435, 51.767671285513615, 56.68567520993454, 61.45047442462325, 64.08782296054973, 65.4070308069372, 64.8908879986994, 64.51357439904598, 63.18474426952027, 70.73530268464715, 73.2966852410989, 75.6403687067986, 81.36444195161162, 86.4288940054278, 90.68463967284606, 93.24660554280234, 96.99889248733841, 100.74530667170635, 108.00409332878169, 110.85411867562179, 113.1605583848586, 113.51399402326078, 117.56838107154871, 120.32201876310504, 125.88657798863377, 130.69300296828385, 134.56878488614183, 137.6784612266234, 142.6332574682997, 155.1945872263281, 175.190631664925, 185.38681366086735, 189.52653578629386, 194.58872275813212, 203.40533561136337, 216.69494633580618, 223.8472408501089, 232.72606667659667, 241.05349307458513, 246.405352710962, 250.54578888915756, 253.7572464253972, 260.8923999002917, 267.71759441370244, 268.7551336843527, 268.0677022814479, 259.44453086302576, 259.0969033913326, 259.6524235667075, 260.0581171338283, 259.8325613906969, 259.1395359980724, 258.91329344000513, NaN, NaN, 24.43792053931263, 23.80777709125267, 24.946446452382716, 24.903353926049622, 26.04214353447002, 26.40830578261529, 26.550991395870632, 27.46810154403357, 28.163333941926094, 28.600386089706113, 29.99275411311118, 32.010472222809895, 32.85083056954774, 34.207817326267985, 35.30598304204411, 36.0347173704008, 38.20013796532208, 41.138304975771646, 43.631453586637654, 46.15891799987956, 48.09975836323097, 51.03298285493268, 54.702905386444236, 58.22420616193747, 61.52385937169523, 63.05837249469914, 65.33118285297068, 68.92395517324653, 72.2213356661853, 74.85870732216354, 80.06401485329256, 83.58397679604468, 85.41045789701583, 87.5322107099179, 90.09907771898546, 93.91484888752154, 99.93546421619266, 103.81817264455503, 105.6549956432929, 105.4975414099163, 100.33184795350495, 97.93819750647187, 101.4350244656608, 106.21744836580389, 113.57001329750972, 117.9904333965592, 122.98494000572634, 123.0212120192288, 125.78761180372912, 134.63218207818124, 146.0710282120277, 166.77523126462168, 184.3598433515052, 196.92297319389723, 204.77260189031549, 214.68401759381848, 222.39016810784926, 231.22337994034555, 239.3032884801615, 244.88335154925892, 252.64001434642103, 258.1584425565788, 267.2184352219339, 272.8759958090688, 268.9699864885049, 259.0284536977178, 257.65829471412434, 257.9596029639594, 258.24087588825086, 258.42627616698826, 257.87987997465814, 257.65900832709667, NaN, NaN, 21.926067469759513, 20.88994495909107, 21.07088911819067, 21.39728843480311, 22.240112300047993, 23.927079484539377, 26.058079612694623, 26.899169108660708, 28.29355276643143, 29.83518409074649, 31.59726278304659, 33.90806363711687, 36.80771071668427, 39.00664966786289, 40.17653952880449, 41.714484677500224, 45.01877133153329, 43.9823317550211, 45.88413590610227, 49.73624464869282, 55.24112545339122, 58.09863077774992, 61.17182636473308, 63.815131993017424, 67.77862707687272, 68.14059994179699, 67.32716976153172, 68.05670498944727, 73.3404626004439, 77.66755357792336, 80.82063535638578, 83.01730848563594, 78.61527571717288, 83.01282574285561, 86.3149019177085, 88.07043387015196, 86.37741464240747, 89.38858658692166, 92.09759645759313, 96.64381176219916, 101.67403069687217, 108.29024118696357, 115.82341197860566, 114.56503932743165, 106.87999098545674, 110.56559467362263, 115.34953743119162, 125.1165744162423, 140.21508650426597, 161.09578847866757, 177.60652818755182, 191.53234711356416, 201.4331748544141, 217.56062705534328, 227.30624042067666, 234.14341576363455, 242.62774394458987, 247.94698726001465, 252.55306435472846, 256.9794211380594, 263.01765852964195, 271.33108189979504, 264.3779153146528, 257.4145536225233, 257.1499971839406, 257.3654798022765, 257.2179761848905, 257.1121214227533, NaN, NaN, 24.24587341855864, 23.689793735006983, 24.6073400007011, 25.301411560183034, 25.77504870038823, 26.2113143855191, 27.7162605635319, 29.146950322001587, 30.097709636089938, 30.129017937481247, 31.710009977113575, 35.20348698851643, 37.95965571898733, 40.640510781512596, 42.28729513571201, 44.48695195636518, 45.66116394203341, 45.3618216997713, 48.74102765563252, 52.96420490014371, 56.78125567816975, 57.95981477011951, 56.345477631235376, 57.44370558024009, 59.786544129343675, 64.11657097788014, 71.38558977714311, 73.44588456695186, 70.87275862934563, 68.22255635823626, 69.0963119573069, 71.87623739724636, 74.95226967077046, 78.46294956319757, 80.8741045163607, 85.64209627483494, 89.38041814898756, 91.65396010786961, 91.72807135033568, 92.15750427066163, 95.78645685234783, 101.53693724709221, 104.91433350407428, 108.2970538252973, 105.67160975707223, 105.97664575074892, 110.11077640790987, 115.29316843913716, 122.37735464368713, 136.68933046467413, 150.99335246713215, 162.51001880100185, 176.45055481772093, 191.87569112034723, 200.92356674347536, 208.88713993826434, 216.09981729618775, 228.02789895538297, 238.19408151848393, 245.92236599871913, 251.38660706986735, 255.80758927737878, 263.5785615057948, 271.9652875344312, 262.40818234327025, 257.91531521303654, 257.57824611083146, 256.6986718727221, 255.8112827774888, 253.1192690254841, 251.88834131122002, NaN, NaN, 28.646167822279974, 26.099265175847286, 24.768485261756485, 23.58696910484386, 24.099647198496324, 24.68518159280128, 24.68028804041213, 26.332611140087526, 28.723151028290655, 29.749527359538323, 32.47209474472288, 35.85738996187272, 38.3554713666773, 40.22433236756791, 42.611143197545296, 44.44762730976556, 46.24219034315523, 47.88433381668984, 50.375381609393415, 52.575721741815656, 53.931498430907524, 57.15952353220539, 60.23623691678691, 61.33289882976706, 65.06602258378433, 68.1381623293811, 67.10112810588812, 66.79762880598852, 65.68777156646146, 65.46191589992331, 67.9508850091357, 74.0353039979124, 79.9076825069974, 80.56966965523593, 84.16837112217728, 82.47880130024157, 85.11538913508883, 88.6321934822163, 93.10073429611343, 97.64117475238774, 99.91416569638515, 102.11538088984223, 106.3486059372407, 111.11688915750793, 116.81718838904722, 123.44754058615231, 117.98821992387224, 118.75186472296559, 138.42231414533995, 141.96001141940636, 153.6303236133902, 172.02109810041736, 187.0183026610497, 197.9557428482817, 206.65804237209576, 217.8455136466212, 226.86145908501157, 236.94121967154337, 246.20538781512698, 253.84775640047724, 260.9418237879431, 269.53774081689517, 276.5799189004981, 266.1597598359126, 257.2112764435181, 254.42338388157887, 253.59244667088734, 251.7619976621675, 251.19407890065705, 251.1620731251481, NaN, NaN, 26.515499840422287, 24.963093943617356, 24.592024630105392, 24.147145774093794, 25.10039901062726, 27.748811020495513, 30.91139236454966, 32.59913979667602, 33.476084330981124, 34.499733652809894, 36.26517943076946, 39.86540512092128, 42.87830040881269, 44.93339391583883, 48.385625150695546, 50.07048225757921, 49.92153570133954, 54.548991235151114, 57.48304762962207, 60.34356040762713, 61.69299521865659, 63.44826077093489, 67.11099221409509, 70.03496600626308, 72.378647144374, 72.8850164911555, 74.56362537030098, 78.81128801762816, 79.83083755799545, 77.76779663922932, 74.08969471259655, 75.69615710566514, 78.49010758413617, 79.14460165447262, 79.35946728653488, 88.24001861982167, 85.38593841913455, 80.23465218491373, 83.5290002802933, 85.5898399687904, 90.25103905830271, 100.70906201591515, 93.9840748587228, 94.42151662984485, 97.94911238998145, 107.65295685524364, 120.17159336253768, 134.9079094882374, 151.90262643501293, 166.2680506643831, 178.14821855713376, 186.66454454010224, 190.28357374558328, 201.23749006205912, 218.35317245083937, 229.71714386530803, 237.67388299358257, 243.36525278672607, 248.8206822482705, 254.2431026525764, 262.3662636815895, 269.3569349716964, 272.917856122656, 275.86655383886813, 263.36721191546246, 254.79898948989955, 250.74947396480727, 248.76740962093595, 248.73714403176012, 248.69523432053722, 248.77395561355624, NaN, NaN, 24.989584065257407, 24.616037194608563, 25.569927886735865, 25.566042259171486, 25.928327978739212, 26.768989309299087, 27.869808139185515, 29.153771597455727, 30.65893467369035, 31.6837778060008, 33.29949999758359, 34.912465369248714, 36.1583510790379, 37.403463665121805, 39.1978721219084, 42.39080004876836, 44.220856779491, 46.19928026241305, 48.98732862132716, 52.4699963419285, 55.88524973209214, 58.304376209989506, 58.84688931816398, 57.185905139563964, 58.16871809639664, 61.02837415979725, 60.2512524635882, 62.77560369942957, 65.8569177329629, 64.53644709383167, 76.41943443655332, 83.7892337118572, 82.5789108392261, 89.39521111056372, 91.38064162811403, 93.0229439489737, 97.53911450120212, 98.65084596272125, 99.20179900811445, 99.8637067281597, 97.74806513606234, 97.56191600321273, 99.40401727101884, 104.54644822075802, 110.41820233334906, 120.73826043471371, 121.69441772603886, 120.97857995221857, 135.3254222238476, 145.84955567505978, 157.87521643291478, 173.6542485712516, 193.00356528915057, 205.4581506965573, 210.73497560219448, 223.48327039199197, 235.3193343597199, 246.14785992257657, 252.63230841934043, 258.4190999959321, 265.4371718402254, 272.1936235239555, 274.1950208539454, 256.4367242864153, 247.88863478216385, 246.40535392946762, 246.3821153081512, 246.71231115083714, 246.85442455078208, NaN, NaN, 25.66189851325594, 25.734814427889496, 26.39367286243504, 27.750579806164485, 28.446026406416824, 29.213183188239327, 30.459911395621592, 31.409140628777656, 32.912209722333436, 34.56526408405398, 36.071185145060824, 36.950111698724534, 37.3515539713962, 39.51502243772214, 41.64427180101646, 43.11088598949343, 44.757762678199214, 46.11250948123013, 47.872202445209204, 50.694480721723394, 53.44718499478046, 54.90802312766749, 54.167458734499085, 53.790635672521034, 55.02739567880221, 58.99182828670009, 64.27871024495452, 66.4745168300899, 68.67942747986429, 68.52776177979082, 68.89336428867928, 72.11802174364065, 74.54480670062848, 74.76526960018464, 75.57174392304984, 80.85582901124704, 83.4285005386019, 84.15138966710177, 91.47724165401122, 99.61911132548086, 103.31730832717514, 107.26745510998559, 110.04843977355003, 113.99942534187805, 108.44846989194505, 99.9451240776545, 96.42253556607908, 104.2105145098451, 110.54805784768233, 116.58330828998542, 128.38793206398776, 138.71198929246333, 148.3132186456414, 165.12902288005574, 175.83021417429197, 187.57319386504435, 199.54947195038602, 210.3352701800232, 221.25611467096948, 230.06239478679035, 242.53797484593116, 253.9058345514712, 258.01300984934784, 265.28363698071234, 269.88539029586843, 253.84621217113616, 250.55695693696345, 249.82250246208673, 246.86022451344877, 246.25148256400135, 246.5109504679832, NaN, NaN, 29.690231900562647, 29.244986257575732, 30.86344539971782, 30.932079205059605, 30.813918531066875, 32.7250844476381, 34.598600664762756, 34.4832528140748, 34.99735037826519, 37.64150062303981, 38.480044319580564, 39.284697875381354, 38.985812935705475, 40.26391966290119, 42.025916280161766, 42.38758402032404, 43.487364881452606, 43.11338591699103, 43.62123041263148, 47.50964018808004, 49.86019847587314, 53.31615666740981, 57.0626041878419, 59.48209673680923, 61.67431351500301, 63.35789852481507, 66.15741894086861, 67.76689253785273, 68.71101751623056, 69.72234160856327, 70.68115097602306, 70.60331187053227, 76.02446158662252, 81.95991908614127, 83.49749622066261, 81.29803866265526, 83.04942581493312, 85.62544919747276, 86.65907796062659, 87.98200962705118, 86.47591946332938, 85.74722464571221, 89.99912043126204, 91.45729162170568, 89.98209669480188, 90.85467616319394, 92.90233698445763, 96.12993686544716, 99.36722327779981, 100.10194169262338, 102.3029126295406, 107.15537739430152, 114.37120787917979, 126.45796604113218, 142.41358705817112, 156.60290511255772, 169.6378875475922, 186.11100181481433, 195.02021383759578, 203.35536782458396, 213.8940684230413, 224.6137671911889, 236.05454790567384, 243.7267361513708, 252.2498666911346, 261.90801690686254, 273.96084452353114, 270.31912331724993, 253.77293733042558, 251.077788561907, 247.8192717245169, 246.50999361074986, 246.6130551206084, 247.0344905511482, NaN, NaN, 34.71320096478976, 31.97779457263616, 32.11992568705387, 32.77516198932165, 34.02236844915583, 35.008122818227875, 36.06905602075319, 37.34973457826747, 38.59215141564203, 39.98237536647106, 41.37113994978006, 43.056556730874554, 44.70463679060025, 45.576845926539285, 46.85673355765967, 49.28231194276417, 51.29618559827608, 52.977811780611255, 54.69714237906127, 56.71057512686072, 58.61967685563262, 60.3719887160458, 64.33137936002366, 67.44990575779707, 70.34072943729788, 73.01234921391426, 75.46757405882839, 75.0647621181454, 72.72640317236305, 72.72452337148225, 76.2836987632187, 77.78585499313567, 75.77597157918846, 77.24459670515809, 79.53260023737624, 76.55915866101573, 78.17780131465418, 78.97326683142356, 80.09369213265626, 81.51536184988647, 83.30366172617673, 86.04905182387195, 89.34513498883142, 91.5415593282839, 93.9293129408821, 95.95557475883389, 104.0567607462972, 115.84353524656889, 136.66252853329993, 153.6864216510719, 169.6088191647593, 187.02375496236024, 198.94672870390048, 210.19987620282743, 222.02524360304588, 228.63479912486613, 236.21625568037103, 249.23901658479951, 258.58757427710964, 266.78663647207094, 260.64804268107946, 251.3838021694683, 250.57088973561028, 249.72830256921767, 247.36956715739524, 247.32625876535946, 247.60845015124224, 247.68256429407234, NaN, NaN, 35.04891865401775, 33.60451837412457, 33.781331851759475, 34.25005894409403, 34.82933985125052, 35.70479637077427, 36.652552474220045, 37.71197063307605, 38.76953489817065, 39.97422395463483, 40.95736149281179, 42.310678508227575, 44.51409203274433, 46.89860433903439, 48.35860484239885, 49.6705616003093, 51.4273921076081, 53.36583051152655, 56.08041692583659, 59.38571602284323, 62.31872854643882, 65.03173192675773, 68.63437456703393, 71.49757611860835, 72.30781840180956, 72.8827178838547, 72.22115325826881, 71.39791863056145, 71.53296196076042, 70.73085972088727, 70.36985501583605, 72.06172056146707, 74.26328567002354, 74.99986314945339, 74.62685892767742, 75.27692506588318, 79.45879751287944, 85.2545398980029, 87.9663735757409, 89.49817267159253, 87.9474140164083, 87.93599025364232, 90.35208290867436, 93.64862434495625, 96.0705090977932, 97.6139444525608, 102.67969044937648, 108.85997615643595, 119.69087639937395, 130.5299234700397, 144.2551758698743, 163.56871150238297, 188.9454671580061, 204.787108645491, 217.21263925472056, 230.29609039528626, 240.4976762920033, 246.03144161010107, 261.20660404603706, 271.5501736756411, 259.786134225145, 251.28014409421846, 250.57023154154155, 248.93351880642876, 247.28302292243453, 247.53696057293433, NaN, NaN, 31.832306540247792, 31.311313489063217, 31.7846097384506, 32.18068634529246, 33.02229629827147, 33.713930493800405, 34.776347243561496, 36.02152541144828, 36.93417710815326, 37.84634833833188, 39.05356295551471, 40.22366160211912, 41.72694567372814, 43.33898443234353, 45.06231625599101, 46.67290659331661, 48.06236583631244, 50.265454576108596, 52.1318559553503, 53.741485679985544, 55.79260354399952, 58.32330777295448, 61.14551124276491, 63.37666068942275, 66.56950554185897, 68.75594102512964, 70.83821827524271, 72.87901410168463, 74.96232968923105, 75.34480159705575, 73.30258631079532, 72.89723784883745, 73.45070035479513, 72.79200705118167, 72.24291753108861, 71.94183046279855, 72.71740974520664, 76.47203149332391, 81.0350522622591, 79.93118369975593, 80.87832681916099, 82.15503408376048, 83.43117453885802, 85.07517972397883, 86.71821824529378, 87.80726206802633, 87.79045351593469, 88.50814838534883, 89.77945173844326, 91.24080467214344, 94.17233609624655, 99.32134391473352, 111.48878636979413, 132.90468751374348, 154.1223351660923, 171.8808628001419, 191.577425325138, 205.3346334967696, 215.4331683311615, 223.3909805532357, 233.62671364176327, 242.83095579161994, 253.0462648504284, 258.13514322049383, 265.72209248229296, 262.2528099242281, 248.9916113933234, 247.63491474544944, 248.1759660607555, 248.72097839342766, 248.83310446472876, NaN, NaN, 31.276271965825707, 29.72123751646366, 29.78940682950354, 30.557015273586224, 31.471815484583754, 32.459328722478595, 33.817690590868175, 35.35926957353821, 36.973143536515806, 38.734604032446754, 40.680606274028904, 43.14373559435305, 45.19793107211655, 47.32527365893286, 48.63873065177279, 50.02474203879871, 50.89379881438844, 52.4288945462606, 54.0368866098908, 55.75498420024881, 56.8810699174464, 57.89734465009098, 59.50248330828927, 60.66548647276331, 62.567772043706015, 65.35309883672754, 68.7987147846757, 72.83649140125841, 76.72320551748716, 80.62270096342358, 83.36107954975236, 77.1328091329677, 74.2964059547507, 73.56984200090619, 75.26316166441445, 74.01403175919457, 74.75354588210196, 76.58825845754308, 77.68809937480088, 79.44890553334452, 82.08915621320492, 83.36517491055328, 84.89705879594489, 85.91334674694468, 85.8937359834019, 86.64903656531746, 89.71263960452042, 89.95244281386431, 89.42243022704965, 91.47052271578181, 94.02833852736933, 97.8878077140294, 107.43202581266566, 117.47820617137762, 128.8426065686188, 158.1133865124092, 181.91697724427755, 196.51487852595127, 213.5892931153943, 227.04002787346553, 233.99550789331147, 240.24009993209214, 247.6987230030346, 258.8467882840288, 267.35858686569577, 270.45386387796987, 264.57622942206393, 250.08645148627394, 248.11665872727892, 248.51109904808462, 248.76052608160626, 248.99975899376025, 249.1173786726646, NaN, NaN, 31.018733759957495, 30.202213781188703, 30.639944929151852, 31.888338241708414, 33.02387091108916, 34.49278799489708, 36.03310790176392, 37.240205775890054, 39.03964021758171, 41.35421684924963, 43.37319561917121, 45.42894703054565, 47.78066618525499, 49.609861228697866, 50.331893686569785, 52.27488869146992, 54.1779077187572, 55.711126540945045, 56.72521525634331, 58.25934463316896, 60.23494360683074, 62.6164545157576, 64.62398721549516, 68.14798715897783, 71.59258443123028, 74.10994747823145, 75.52057984977436, 78.2653150966321, 81.7871541032404, 80.06977433343398, 75.51506654080858, 76.80096989123896, 75.9681523366046, 75.53043583474737, 74.46745381162525, 76.53667293021883, 78.04274362832867, 81.24608654975631, 83.04030012171329, 83.90887760212284, 84.96115980296783, 85.53653778155591, 85.8177509255454, 87.86532749827307, 86.67071601649741, 89.0021607515098, 90.1593984970548, 91.02604716710498, 92.76945151900279, 96.87155332214819, 103.34482646832227, 107.14772486198324, 113.91483610135653, 131.64815437105904, 167.4406237582602, 187.31443775028907, 200.40841771852632, 209.6741588594849, 221.66315235329972, 230.09916244371215, 239.33793132060245, 247.78629892506123, 253.78099109585872, 260.65615870546424, 267.57687245903116, 266.49326404502614, 251.24351932628173, 247.83260845889572, 247.77981163294817, 248.1903562055703, NaN, NaN, 31.127543213032414, 30.23950784724656, 31.084878315393805, 31.9256214888052, 32.765706713364004, 33.569024382131246, 34.44379365904353, 35.06009650507363, 36.41656742508945, 38.47413403175684, 40.12381649526146, 41.88436331546095, 43.9035575024549, 45.84906213456533, 48.27201334001976, 50.10362776124222, 51.78687833024598, 53.434614262221146, 55.710225126173306, 58.28065841183645, 61.07084956205043, 64.0419957226361, 67.418149756365, 70.45553429938487, 72.82957514494024, 71.14330453242889, 70.02911694571816, 73.61221810531138, 77.61957602780241, 74.91803795066933, 74.90053915666962, 76.15734152134267, 75.05590264672726, 74.24753869406233, 74.6564912434866, 76.79935340684723, 79.0846554586701, 81.58002783269639, 83.1951466372883, 84.13399212267987, 85.22104761625128, 85.79932689027969, 86.07330808587578, 88.41177419170522, 91.03740472727377, 90.13558823163561, 89.8256806318844, 90.39421283358531, 92.43405338912149, 94.47598016355636, 97.99453769550266, 102.39699886069288, 105.90691223224717, 111.50218307165959, 130.69723463964803, 152.86724264727127, 187.35592721499862, 215.1851090594601, 235.46199412705195, 245.11804419515576, 249.84166537923318, 255.48233180828086, 267.1211666388427, 270.9559531561329, 256.0973229343381, 246.20168949741173, 245.40671024495992, 245.9556363098122, 246.20361971103233, 246.453012308101, NaN, NaN, 31.12576532992435, 30.604097121935347, 31.07737334375531, 31.65896939913146, 32.46286852115787, 33.377005985195225, 34.32666736749133, 35.46147426376436, 36.44807342902628, 37.6193784168242, 38.67881332619459, 39.84971247398233, 41.020726794691335, 42.33840613965933, 43.508597860920716, 45.194794599042936, 46.99100421421842, 48.637760833418895, 50.02647530215452, 51.488675360067035, 52.9150456851118, 56.66816647097781, 59.749832761379515, 61.47099217450814, 64.12234026512246, 66.07232441511465, 68.01779605894859, 69.44689968697958, 70.04594146332518, 71.12200694584413, 71.2322508227091, 70.23303623449635, 69.45794903308935, 73.69296413116095, 76.6246631250463, 76.77033482846221, 75.17093051992569, 75.48945880356375, 78.50073634092696, 79.42032270685647, 80.30768372117812, 81.39717842299099, 82.4842214323531, 83.5714097684404, 84.43929536244318, 85.75351540201845, 85.95950433614212, 86.60658915062832, 87.91754064119625, 89.2301615359108, 90.09677584065322, 91.40326332190615, 94.25616896606434, 99.76854337105391, 105.27309722935267, 109.23436582659126, 117.85138281098699, 135.80003476294254, 154.8632065585075, 179.55491621044584, 198.19504874623632, 214.45396842756927, 226.8744270061918, 239.7270554342664, 243.80810503226002, 251.67844603177483, 259.56171475124336, 267.38405077008184, 270.01231972322176, 254.15259378530035, 245.89157392780805, 245.6920638906471, 246.08540824915082, 246.49338482005948, 246.611212370421, NaN, NaN, 30.572713798211957, 30.051369150168316, 30.34050526577461, 31.07015868431444, 32.058660396476554, 32.97121807244155, 33.95753265515275, 34.83257285606007, 35.85440888764538, 36.9120193981266, 38.08093581828386, 39.24871619234788, 40.454415938814435, 42.139170247083534, 43.89754807758341, 45.72754012022429, 47.378553517180094, 49.395060506449205, 51.0788153201536, 53.28087544565859, 55.667802589545246, 57.64868224572569, 61.20823654778519, 65.03397772215425, 68.41306604232429, 72.27619628459894, 75.32019360302688, 76.74568077275107, 76.71183028809472, 76.04820404524436, 77.47664792328148, 77.69362602710378, 74.76020809868217, 73.9530929667708, 75.26366338390912, 75.5138607432657, 78.92569897945566, 79.43899699740335, 80.3935411340752, 82.96101245509362, 86.0410993490456, 87.68246626126395, 89.13565343060716, 90.58804242359687, 90.75690393036881, 90.74374199854432, 92.75305330729634, 99.91601815630622, 108.18860690786337, 115.1792117565081, 126.23788943978536, 144.49908590766904, 161.4693934282793, 176.2670512563075, 191.9362031285184, 212.88538510062185, 229.88965837983713, 239.89348643412418, 246.740139295779, 252.0713958254387, 258.52063477204166, 266.9303538143912, 264.37210100145046, 250.28484342926316, 247.76324248353927, 248.03426422354195, 248.30560834972235, 248.43907974741558, 248.28055828114225, NaN, NaN, 32.30349550980775, 30.712948324182495, 30.965243823581428, 31.9912138326274, 33.05426929262353, 34.18997537895971, 35.28857262744006, 36.793569611156514, 37.81663887338937, 38.83800486152694, 39.97152311991593, 41.06796831196271, 42.23735988970897, 43.073226264344726, 44.57641325695346, 46.4097899283729, 48.13172039566214, 49.59592085583692, 48.90033704785204, 47.68109734577815, 48.62820976814826, 51.858623913590506, 55.3068236850194, 58.46912818798249, 59.78494652287947, 61.983660181646385, 66.09696464587464, 71.75303923259008, 76.08288139230893, 75.49408687648354, 77.99835576368224, 79.39371934916139, 77.40319080664251, 78.93793568217956, 81.87006239658317, 83.49045523339208, 79.53432370344485, 75.1251794166773, 76.44922146698359, 78.34850010715701, 80.36003310387073, 82.40500277811385, 86.80466599453769, 91.20857896666863, 90.76953121382455, 90.61342978127833, 93.69787058244104, 98.25255682421377, 101.04126211969145, 104.72461306992709, 112.23705582289352, 124.16659406204711, 140.51888997531498, 158.13251108224307, 174.12460816643338, 187.51568295379724, 199.3945744229269, 210.2401642825473, 217.6219658538913, 228.87354733571482, 240.43720316664087, 249.0607199920078, 255.6650768140921, 262.20489001244687, 271.1403706276548, 262.71421785024523, 253.22740097834807, 251.9818847274449, 250.32447990749725, 249.3370125702319, 249.52237267704567, 249.7186946502589, NaN, NaN, 31.453878870158313, 29.93662756974344, 30.374015944811575, 30.88106397556543, 31.978182859493494, 33.297148364104224, 34.948832946439005, 36.084436073485506, 36.739114153934544, 37.46889861266713, 38.20202492168333, 36.57778246453337, 36.78917198887938, 37.26259895355948, 40.273811993763736, 42.442844520397045, 43.83531864293091, 46.44196414976077, 49.818717019666614, 52.86928600052106, 55.4369129270146, 57.70673334732609, 60.64190673250377, 63.14273905929381, 65.19927370132531, 66.6640725129415, 69.08553213542564, 70.76432810116036, 71.42596841783997, 74.9409050787504, 77.72980966533528, 78.52902626253055, 81.1638154790051, 81.8222285981796, 83.64521749547052, 84.59587827217132, 84.95363407936814, 94.05177787648209, 99.11670648514846, 101.03102900371545, 94.62006307990133, 87.2841472319257, 87.43046320407409, 89.92258608287754, 90.35531336610227, 93.29102383535772, 97.84859468123483, 102.27042985625536, 108.4500882051216, 123.02984768529491, 136.00483072803084, 147.52089734062952, 160.3984185158366, 169.42814048247675, 186.46902176153952, 201.96967964316056, 213.81857558950875, 224.50664880335697, 234.33118841531464, 241.56386407896582, 248.28981103340345, 251.73566014017086, 258.1199513423866, 263.8995490468864, 268.79143966315877, 270.59940554977163, 259.45353066170185, 254.73191667701158, 252.57380546893933, 252.13296881911825, 252.19238586440432, 252.4846446865306, NaN, NaN, 27.768812430308113, 27.765099670948647, 28.574366796829693, 30.189475493046864, 31.547833004689128, 31.874550279686147, 32.30821549173103, 33.185589900496836, 34.83580696315622, 36.59448136021741, 38.60914382961361, 38.489504145886876, 39.88107264847384, 41.70964894789295, 42.21545519577696, 42.983522483563775, 45.44050846320125, 47.124555510659796, 48.84604527224133, 52.185738858988145, 53.976699583497606, 54.410922640332274, 53.5191315365532, 53.72824422364281, 56.477214107101446, 60.544785435638694, 62.85814336862676, 64.83796618795263, 69.56673483777261, 72.87006561809709, 78.25583509554474, 91.02219671456967, 98.82742282387369, 104.99644466634669, 105.87703704260511, 103.78321390808392, 100.47587938741187, 95.64402464495639, 87.83294469907833, 82.75967353842923, 85.90190919523903, 97.4951416006314, 108.81609771341849, 114.39613576852898, 115.441396887559, 117.96245409938771, 115.04638316838752, 119.33602602000029, 132.47258166358077, 141.79775725212355, 149.76632330212124, 160.26155176933997, 171.51537172270127, 187.6769178972327, 197.05093436682344, 210.0868052340431, 221.20155508185678, 229.19620991142656, 236.5499197481025, 242.99978971862754, 252.84007294540206, 261.398202904675, 265.1425382354508, 264.34145049101033, 260.42618465225723, 258.07981107633645, 253.6394349132274, 251.3163022328276, 251.19615788009565, 251.38869596420292, NaN, NaN, 26.90554268379462, 26.496490604059233, 27.082594831377424, 28.40480368034496, 29.615968146326182, 30.64338794464205, 31.262290815350003, 31.700882105526308, 32.393330877613145, 32.90349664323519, 33.63139570344076, 34.58178037799125, 36.19534605375444, 37.66143612487096, 39.79013890895484, 41.55162289557492, 42.024256834145795, 42.60919283366999, 44.55116476107108, 46.97035671922825, 47.84424799822285, 48.20745898978929, 50.484105609815245, 50.99543526913046, 51.50549255015251, 52.82526824408775, 56.131438897712734, 58.698377228715, 59.430210138667725, 59.63954044940738, 61.9080581179881, 64.6968156983171, 67.8477545654906, 72.17123973498292, 78.91648281515555, 82.06257188192848, 83.59584903856292, 86.97765082206979, 88.14918760913785, 88.65363263142666, 90.55349417340466, 91.14867363804541, 96.57082881715694, 100.97384285272969, 99.37382054118477, 107.58783129590465, 116.39602564237447, 125.35580440277982, 127.56228228333758, 128.05970617855078, 126.49517758484589, 131.51040918734734, 142.9726123944833, 154.0249916699116, 162.25068280643725, 173.51590009196073, 187.02787274827105, 202.3643873731648, 211.21578351493505, 220.719947077897, 231.57660341127277, 241.44537982425777, 252.41471139287248, 258.76179294492704, 264.2653487713598, 258.79514746483426, 257.8419155913624, 259.235843356064, 254.86173767596728, 251.51093346954573, 251.13489660052645, 251.33052504275997, NaN, NaN, 22.590633520711535, 22.73542585409346, 23.654653807871473, 24.867069309021016, 25.785013171521122, 26.812810285355344, 27.802632811159363, 28.606982251500245, 29.227543427805976, 30.18101023821369, 31.17112353226026, 33.9258111663972, 36.45632662395787, 37.47968958356829, 40.08810426870896, 41.335945333846226, 42.17770595980678, 43.38229066374998, 44.62640410254141, 46.02351198309061, 47.52975244356861, 49.22355483656848, 50.61441547235652, 53.18329896805921, 54.13094972906463, 54.857675705573726, 58.00873915349203, 63.72953148017463, 69.15577135218929, 72.67629107282815, 79.05928829549198, 85.6575312179935, 88.67083188751963, 89.83516474601899, 91.44951842383782, 92.70767215407378, 91.97260097909196, 96.36795736074872, 97.83368836283037, 98.0506199469325, 92.9656071795923, 102.7075939559894, 115.75866095177888, 119.63069792652703, 133.5935437897833, 137.70547452122563, 144.58718430231045, 150.3279050986988, 160.32560680588398, 179.81916734683068, 192.02294875327848, 200.08792409442938, 211.8503916217387, 219.42361529116016, 228.6237952312673, 237.52261000674213, 245.9763708588244, 250.7694307811263, 257.1231180333246, 263.0331518001138, 265.05235341346656, 260.6091613445225, 260.6323635997416, 262.1057291517562, 259.0077252466318, 250.88028560459082, 249.87042208430498, 250.0356585333571, 250.23336380400144, NaN, NaN, 24.763353866852533, 24.39053816243908, 24.607442622487625, 23.055486869129588, 22.717966208047525, 24.220549024787665, 27.013969887233852, 27.341744920383995, 28.62339161825995, 31.194871538025115, 33.69141302766181, 34.38345689910105, 35.44384552984051, 36.46898748985221, 38.67283962754567, 39.36326597823664, 41.23069335414185, 44.89965021173144, 46.988936851281636, 48.78306793267578, 50.542990237994246, 50.02026679537336, 51.03965406478158, 51.98542292548676, 51.83355868399242, 53.8831196478091, 53.58423386425715, 53.87638300350358, 55.49130677992174, 57.25128321864985, 58.34872308541709, 61.42307107957202, 65.82493951832078, 67.1371610166386, 71.45681606690829, 76.21950605053863, 79.21805397592509, 82.57895260060036, 83.59613333214051, 85.13468275755541, 88.1841037771382, 90.38614976077636, 91.11339905022973, 91.83653504089214, 92.38783520606748, 93.49253940032513, 95.89378669965329, 97.54393151442106, 101.03095177194695, 106.54909925503708, 105.82867392036056, 110.24944793440113, 118.73415410217163, 126.66422065976917, 140.69006874946072, 161.33710586562657, 182.64786068118596, 195.54013560221279, 206.41070571883867, 214.88662535921904, 227.9243524064476, 237.8494343540582, 247.92636271395182, 253.21690503783893, 256.52282600930357, 262.8124759157928, 263.474486815852, 259.8170566584943, 259.4016611699454, 256.89780163031287, 251.75237251627564, 250.6175280037892, 250.6671310637535, 250.86081484213082, NaN, NaN, 26.82709910476046, 26.34443878816549, 26.780991383527052, 26.371099922526323, 23.456764546998322, 22.60462120157383, 24.551502406749307, 28.19136710582883, 30.356960345425914, 31.787153152424132, 33.624374206472034, 37.1867700101046, 38.280943104629166, 38.38270840182804, 42.01400855220372, 46.196008300418285, 46.9630594689357, 49.823774432652286, 53.5301631443636, 55.84177073104801, 57.780615216634644, 60.12219268734166, 59.89493649346101, 59.590563568734886, 59.50583296797319, 62.219557355089655, 66.54552389510391, 70.43031279614259, 69.24610971060234, 70.19256080066953, 70.56320316999089, 72.10564204417034, 74.96570519340312, 77.81855523477127, 84.85276252126977, 87.84816139102739, 90.70022108393097, 94.58316477351924, 98.9127732425583, 98.550414180358, 101.82415157134731, 95.42371147153942, 95.43797802647502, 101.0894170772426, 102.64136393330627, 105.73088296642905, 107.52296248676963, 109.08252806211908, 115.02427793056646, 130.23010494476324, 160.8837302161706, 172.2323924279962, 176.394518682924, 185.01162799244267, 189.322746345808, 198.21845535555468, 210.79795711382778, 228.23186680070359, 241.9439695821673, 249.10448483335298, 252.99693068676314, 256.0343790967403, 258.78413010057403, 263.28611920146653, 259.9098180876513, 254.5988571947108, 254.22890248495838, 251.9527236862179, 251.8333045810369, NaN, NaN, 19.44532456032457, 18.743181543452284, 19.108577996107154, 20.686918772709866, 22.340589726907858, 22.485068539631854, 23.767966361906986, 25.490986427016008, 26.810615525755463, 27.655178308337018, 29.640254964125337, 31.660002520461518, 33.936134238381925, 36.35854518053814, 37.747416140286944, 38.03835674279269, 40.493145549242165, 43.461982856068666, 45.47882930294682, 48.70440675947848, 48.22390049879022, 48.58279922262324, 51.95836326454511, 55.77514624839024, 60.76045780867261, 64.20383306587146, 70.36344394818322, 74.4702003184032, 75.64050452755401, 76.65879457224054, 78.55834792669265, 84.27586621389196, 88.67729346839415, 92.34247186734197, 94.08851183155313, 95.25402060018386, 96.62499389847605, 97.78529231991251, 100.42054182939216, 104.96719257829473, 110.54397214952512, 115.68272099590163, 117.17255421506027, 111.29734807329005, 115.69645651497673, 118.65244199998136, 122.3557316278689, 135.1966833537522, 143.86163463898401, 156.02916631173798, 163.58360764719757, 164.60385098471832, 165.11167028118467, 173.11944279430054, 195.35156625870337, 209.33328245985757, 221.64275250796453, 233.43640308031314, 244.51135154781716, 250.49230905441252, 253.90491855863007, 258.8592642094928, 261.08470743285466, 259.86827854377225, 257.7121148588269, 256.5529975530985, 255.7315881974956, 255.36007817727892, 254.50561459810706, 254.56127841332514, 254.38941414499217, NaN, NaN, 22.106101399227782, 21.44096061688191, 22.101735847074263, 23.203874914075342, 24.232492381508788, 25.9947223261844, 27.534745202766793, 28.853006735197663, 30.024824572953765, 31.7162883193937, 33.32998021330949, 35.161504318053886, 37.437224097896056, 39.123121394475355, 41.47412977630181, 45.587238488346145, 50.43512820488217, 51.018939331707124, 51.60068577575673, 53.21236971975557, 56.33124177951103, 59.18915091023296, 62.3433719948476, 66.01183842019978, 65.9354961985688, 67.39196927976005, 66.58140795044896, 63.42111977163476, 69.8008071532046, 77.12715030609633, 81.8876030665255, 87.68401818982912, 91.48514611622898, 92.7304013818165, 92.35493311037166, 99.83450860204462, 105.03064814913898, 110.59840628102535, 114.32860432407584, 117.98588722111884, 121.120782115013, 124.06464900591605, 123.90635951902486, 124.66364034401003, 127.97325842937938, 129.82521233395659, 136.4586567742095, 135.0411505279363, 151.26475802207503, 173.44213682970738, 186.45398470480302, 193.7385971677213, 201.43391659429867, 208.21345426021358, 220.27295424651058, 227.5276371643861, 243.01518710899984, 248.01710488235034, 246.39324053842208, 253.8756790482025, 254.9333648296265, 252.60355710812553, 250.73115126311015, 250.633237608988, 248.34547584047644, 244.94705773849944, 244.21502703694532, 244.32631731801354, NaN, NaN, 22.9208058721254, 22.070340754511136, 22.656631039388245, 23.609871561534177, 24.156588212453563, 24.666371045775854, 25.875607186820243, 27.231930514623457, 28.91808448292246, 29.75917710504981, 30.15827630471227, 30.926599980260978, 32.31987577126668, 33.48848805340606, 35.65092737247029, 38.43632760749894, 38.39560842781247, 41.47150092924449, 43.887035333924935, 45.68029006839763, 46.92686559961388, 48.79300931192712, 51.97639117422522, 55.82516996937969, 58.90681243371668, 60.77977916966174, 63.200729630454205, 65.38755317517901, 66.80762981014806, 70.21068668459765, 72.40540282103157, 72.28709150592817, 82.18108792880142, 87.46234493869099, 92.41371793251044, 97.46993048346702, 98.33967779140885, 94.70756111778874, 102.83832252323602, 106.57630734500948, 109.39650514522573, 115.06850846214226, 118.02399822605858, 116.0065803334163, 110.73034631803226, 112.9474191631727, 121.20056689819243, 119.2145818511041, 133.3989300072793, 139.3196657094799, 155.38501166550785, 157.87285672773407, 178.14602324340632, 187.2821858090337, 192.99856199735257, 204.75306201416436, 209.63321185911485, 222.22223400840232, 238.69502319911192, 247.67894832998218, 252.33274598892015, 257.22082142494975, 256.1731926885426, 251.98376191813864, 248.70097903314914, 244.4568686384885, 242.74456939143943, 242.4213774776414, 242.76066240267045, NaN, NaN, 20.885411455232134, 20.586750185256893, 20.95163780157864, 21.648259563787587, 22.381799790513405, 24.035393357891593, 25.13486286579853, 25.608429029560714, 26.70549182152774, 28.060827067870864, 29.085309022666443, 31.24934999330446, 31.541083883882546, 31.86869161594455, 32.41703435727916, 33.919974878061375, 34.9824260397204, 36.95986003317616, 39.45081303261494, 41.5723238055532, 44.50551443823196, 44.793446843499, 48.09383772613309, 51.98338453187489, 58.4381085919535, 61.59080041547441, 63.78379198843915, 64.14450052512002, 65.39331112191836, 69.05658602821495, 72.20356132334923, 73.14453788401808, 73.5749256576735, 74.09112858583549, 76.28579869235816, 80.74657210292185, 83.30506453364097, 85.6477579549279, 88.36163600277884, 88.71894407120621, 99.52490672869428, 121.95801053598983, 119.11168998547512, 103.0765607157291, 126.39459234696322, 134.98051781057057, 134.08627773343338, 130.12874518207462, 132.79689971245267, 142.30511205220222, 155.80008457731864, 164.44617654941456, 169.5622912375288, 173.49795076239096, 177.1951138819147, 187.26718035350086, 200.42642921874403, 210.03689531573187, 220.93006074949122, 234.70741792852436, 249.64541900152935, 261.3752549719678, 267.016776372368, 255.94572366495757, 243.77072125564334, 240.6529913286736, 240.84420337974444, 241.25282820921723, 241.42540259857964, 241.71737522362386, 241.79883226573907, NaN, NaN, 24.870191909451776, 21.548985751910198, 21.398233969579827, 21.39248340477037, 21.756700706096343, 22.340407241927885, 23.810023649737758, 23.880721447269256, 24.61068738677795, 25.56307337679349, 26.809754732581556, 28.423816944531243, 30.402595522007093, 35.03128862426699, 37.30569639875517, 38.843148250048934, 39.34906063279765, 40.589764841280285, 42.34967085931902, 44.694685609679404, 44.87398576617378, 45.74867024685009, 47.17603955791949, 48.49019042883958, 49.368657611326036, 51.122970014427786, 56.07025261050269, 59.14472624337451, 63.20782811324291, 74.53731812441013, 76.73412425623685, 74.96789949696966, 76.50414333407824, 69.12973837308307, 68.13013311268355, 70.43317463071743, 73.5093704765201, 76.03011460997087, 82.06734404297059, 86.67841323385021, 86.37626282756929, 88.57346193563342, 106.15794177857873, 132.98006277466658, 133.64120880860875, 119.58341134480425, 117.39734448742567, 120.48357353809936, 120.93344624887065, 121.16617291822803, 126.46491530723878, 135.7378742898749, 140.36381438352353, 145.2242901995842, 152.08706690299806, 159.62785650678106, 165.83043960218978, 170.72072917874263, 176.11016379977934, 179.1166228524456, 180.38160391766073, 186.7655541040849, 193.33985641143477, 199.70538763967625, 207.47429499973046, 216.29414065778548, 230.64202470607373, 241.54832248085947, 255.18388880766892, 261.56969214803223, 259.00066216782284, 249.65400747483224, 240.96807137396678, 240.62086263247892, 240.88256639597793, 241.28928183744696, 241.4041405835074, 241.51890421176165, NaN, NaN, 21.07596081666763, 22.031135042717946, 22.91175126482719, 23.27268599712151, 25.03309360460004, 26.867716652771545, 28.921702437814787, 31.564222897987182, 36.9258605750022, 40.29986784232019, 42.281462523814554, 43.96483276880686, 48.07172752053513, 51.442397945817135, 53.0472313062212, 53.997191700397615, 55.82196774653096, 58.01528354052279, 61.97434541520143, 65.56712080312316, 69.75049668403062, 77.02076239159464, 79.65989278561186, 73.48995805340995, 72.8105186109271, 70.82270980945017, 62.44689002852135, 63.53752708311808, 67.92862518371433, 73.20415521160143, 75.83586210260295, 77.58597770078958, 82.63919470218532, 106.38410712314817, 113.21786103837155, 114.53044466027556, 116.05144187103312, 113.19282607537436, 114.30819488077816, 117.83464345166142, 118.49630336226568, 117.17733408550875, 118.04668267550474, 121.9982951534326, 131.12628747201904, 138.1851408860533, 144.8019666857926, 151.74442209134352, 161.6707397126966, 169.3686345064793, 174.6746867606108, 176.57880540112387, 183.55247964048203, 194.73135399022848, 199.30991138140496, 214.4851538111389, 229.67679985136104, 241.68314832117608, 249.9250495642137, 259.5485741145608, 248.1228893336094, 239.03664106720566, 237.50540220124014, 237.79338893585108, 238.3105119697117, 238.7235598135505, 238.80927474057336, NaN, NaN, 27.962102287372293, 27.369052051530645, 29.17064482383471, 30.53220987365476, 33.17951843151062, 34.86708799533282, 36.03729560391598, 36.73070240820985, 35.32361909649478, 33.629232732308495, 33.84233974372174, 36.70702424285755, 38.68834444094768, 40.74249009988774, 41.362649988016884, 43.15753400074281, 44.40145360584074, 46.009597637842774, 48.54131050462536, 52.686587804662494, 60.46704352157692, 67.80274577722348, 74.40549520991831, 68.34779535406349, 60.99928902819538, 60.98966348276595, 65.7551908928542, 68.49250069825034, 71.23507240757058, 75.26251265064485, 95.62381327213477, 103.8831328954947, 104.42578680277305, 105.69898334591068, 105.51017337146008, 106.96687518307024, 108.41687950394324, 110.05470921350914, 111.1527183996052, 114.09030528668976, 117.86809624858256, 120.04878580759043, 120.32858058243214, 118.41934890165392, 121.92779681446038, 126.6391055515411, 132.6796586723207, 138.41166832131128, 143.8597757358648, 151.70984367627497, 160.59042421556146, 169.18768596758835, 172.7939137032187, 172.41936380816082, 169.28483876380548, 177.1322464928569, 190.49890253818393, 195.89300982340905, 210.64048673509285, 220.0475275791803, 228.0570975543665, 237.67689389100948, 251.1225805966286, 241.95373094971507, 238.24954948019771, 238.98023240973978, 239.62026347353066, 239.81856024283616, 239.3746885605496, 239.31941670536915, 239.51007987441065, NaN, NaN, 24.830252967193392, 25.047392351841786, 26.703414535800874, 29.12781322007836, 30.337627641151048, 30.772265275225166, 30.766295748703026, 30.758838836213336, 31.414786599927822, 31.960451565588034, 34.494789202989956, 36.804312090129464, 37.90019679850886, 38.88430094109263, 42.95620770868442, 48.12842254566704, 48.23438988499787, 48.11804708450385, 51.19780609750183, 61.21442793208038, 67.78251147997746, 72.73550214308996, 67.22995273075158, 58.96589546961889, 58.40880231997779, 62.98911126344943, 82.26150898501922, 100.43143380064198, 102.99310513028608, 97.47219080722239, 102.24024952209558, 109.9220191242634, 110.62978724345668, 106.95164479634882, 105.66577617942573, 107.11899031760785, 107.84347407978512, 108.91549720879426, 110.91364049488254, 111.81685337684874, 114.33734104132218, 117.08737235118588, 117.81409714058421, 118.19853662483916, 123.70756073139907, 127.55364216711737, 135.82644001049243, 142.28045454936156, 153.0011900262197, 162.99145510550275, 168.82373983301682, 165.46637466459583, 176.22465306212254, 184.24258356920063, 197.7561681391427, 205.9694826585596, 210.93339373115793, 220.97722474885023, 240.2773051444796, 258.327106567309, 255.93536964341817, 240.0725249625431, 239.12315044551403, 239.6722943302141, 240.07803633243063, 240.47937025408427, 240.57912101601434, 240.8392645046021, NaN, NaN, 23.7212444965102, 23.275836837872077, 24.23024921760543, 26.06662998804435, 26.870766979481825, 27.23240883704423, 27.447556163279668, 28.102606690297975, 30.082073678309285, 31.032910060826417, 31.761992725240475, 33.962805785812805, 35.94064899017769, 36.00755377664436, 36.95491518499559, 40.913334176002486, 45.762324159090596, 49.72197213115177, 58.381006185591524, 63.145118423547586, 65.9985591018252, 68.04931038041094, 67.01384742566736, 59.55870412280451, 53.896195929940745, 53.883079071416034, 61.32941939701367, 93.41751022094337, 96.75321343476486, 92.63624068807786, 92.11900531093863, 91.5947714645571, 102.61993480341272, 113.39671055497188, 116.47545555848447, 114.67068106197688, 103.88952292337932, 99.24877137156079, 99.49773982224588, 100.25219132043088, 102.71361971088253, 109.20358433980778, 113.92946722001527, 114.5897161090488, 115.38173245782181, 118.81273821060839, 122.5625000610841, 130.50953256189783, 141.00050206109483, 149.62889135960893, 157.59968193762896, 161.4323882728487, 155.69756164150073, 157.84870374368438, 169.48873995076656, 183.26933841749164, 194.7888397304507, 201.12899765347893, 212.70967806961735, 223.73994532558723, 235.80208355100063, 239.5971268937174, 252.466948844899, 250.41138069362, 239.45085576727192, 239.28913906604765, 239.91643508127376, 240.3219303054802, 240.73731885951065, 241.13844086909938, 241.21672329758334, NaN, NaN, 23.60407283655086, 23.196075167284544, 23.303693803198005, 23.593580917013046, 23.918599294894687, 24.575034959557804, 24.901307039813286, 25.15413190942226, 26.87850153828872, 28.199203234919544, 29.51835898379314, 30.689122337723866, 32.1553746312368, 33.47344684907415, 33.724587416598034, 33.71793605708748, 35.03547309238935, 37.568375531591606, 38.66374497233738, 41.37459281086501, 47.64854061660254, 48.16340605143212, 44.81964995178791, 44.81366418034831, 47.88821495630661, 49.94036947452333, 49.67700159423739, 51.2122513006505, 55.82727457868051, 85.35235901219262, 93.31328149009154, 91.77974127358489, 87.16053342521414, 98.70817333892386, 111.78994948759258, 120.25169104699722, 122.02937711344879, 118.18208067026417, 110.21794760836255, 102.76874192369675, 101.76620658389288, 120.22716342421289, 127.11557402832126, 118.76496419859762, 114.95152820460723, 115.2571517996377, 115.11434096256596, 116.31105656936312, 121.89775298106628, 131.30001308768422, 135.722063410193, 140.44905063196677, 148.10261829699877, 154.74203768188056, 155.16176326904315, 148.92872410909038, 150.88571475704686, 165.36338836659428, 180.37915009982765, 186.66911171441075, 189.5140506942759, 197.453361104683, 208.67090069696323, 218.12061561664487, 225.1829731852108, 234.054586409254, 250.05722506890964, 261.7083568001436, 255.07630349248223, 243.5347370153074, 241.25001835928063, 239.69082111476874, 239.49888094989691, 239.61053160735463, 239.86803832662784, 239.7058221759343, NaN, NaN, 24.4580109062182, 23.570597396067548, 24.600536703992827, 27.3221975021911, 28.49363837584724, 29.298627299018666, 29.80887133690081, 32.23433591299764, 33.11365141064606, 34.286374674747165, 36.56311848468409, 38.10160985881948, 41.25590524563428, 44.19149543265364, 44.55025985341982, 48.21821762025672, 54.01897889583556, 61.80289924113474, 63.63513100989605, 55.62967976812883, 52.60764098835635, 54.951817582853444, 55.67836966167176, 58.16382684405041, 63.297738837346955, 74.89084123581601, 88.8268337204538, 102.17422704065002, 103.19852493691761, 102.17743029363379, 104.66043338708728, 101.42814486912101, 101.99406017925776, 103.16364810246121, 104.18408591118673, 107.11030049741969, 109.73220542232657, 113.11747289623084, 114.86337989034011, 115.43912316186348, 115.95390775100041, 118.88270225944179, 126.24751290893923, 131.53768738206142, 135.94797830039624, 144.2243316972018, 154.40930418519946, 160.77871101846966, 163.6616549202095, 157.6013175398977, 172.2112928971652, 182.3516037259457, 189.42533557597005, 197.44556434857574, 202.94577779168503, 211.76212098685363, 220.62610639564377, 229.89341216258612, 245.01364163532872, 260.95968918141637, 266.61895309938876, 264.3417463833719, 249.3184110487076, 243.21654969781918, 240.44421802571154, 239.68863939493986, 239.37589363504958, 239.08598166966448, NaN, NaN, 22.29020579096745, 21.550649735299604, 22.062886053639254, 22.86791307609673, 24.85051997168827, 26.686540336792266, 28.152678411906887, 30.65066246808288, 31.52752804828914, 32.771699353314894, 34.82419514449177, 36.58480695422386, 38.12126644083806, 39.28988669168901, 40.67885244841293, 48.015340550043724, 48.74655552921662, 47.85848321569345, 48.51435466169729, 51.22575247994758, 52.98611321522519, 55.47354985294622, 58.40694369901025, 65.8904137010684, 67.49683761163645, 66.75331069370907, 69.53910253366892, 74.67033956955969, 74.6614026319757, 73.33309650214521, 79.78248205589504, 86.96694139249442, 98.99275169730048, 108.51711805005111, 114.37506373883544, 119.94486249819457, 134.60457879262887, 131.5348866967679, 135.92793146642094, 131.97467696384314, 125.00073130754186, 125.15300258486816, 129.57863840450597, 137.37673853671294, 143.09669704679513, 148.8442613521075, 156.2377937592816, 163.79870935630257, 169.3812703559907, 165.47075930453715, 170.5778981634883, 186.0215295283307, 198.236979868699, 206.23597343040618, 216.8304771950156, 229.55368489014134, 239.58556872646918, 246.16832880918275, 260.31283384884847, 261.05161092960793, 241.78207102609727, 239.59759015647103, 240.02106951335952, 241.01935517266682, 240.028088383954, 239.38838476840036, NaN, NaN, 22.177805554774288, 20.775623596264854, 20.88243978554118, 22.240288965344924, 23.819171253721194, 24.697909093467374, 25.94425441080409, 28.259230563723598, 30.793540419993867, 32.114492150909854, 33.98516121627875, 34.31130246354167, 35.48244062155612, 37.20470571305011, 39.33224327201136, 40.540610243394234, 41.196115440224006, 43.244663926243035, 45.51879255069339, 48.5620399988088, 50.351572511396334, 52.10776835102763, 55.042669204016384, 58.858096220525795, 61.64377607352995, 64.13271770451654, 67.79937184506942, 71.16720600936901, 69.84374832699683, 67.62959168054552, 70.55371785445017, 69.66981579987802, 74.50340536284882, 76.69651193566948, 75.95590708731022, 76.09305645415114, 77.69888609003333, 92.3484034712462, 93.95429538351739, 93.51563384962691, 99.20355922689158, 104.02644814341967, 99.92308612041288, 98.45786816819457, 106.67059271253834, 109.48732091829439, 114.37375304302505, 120.15688073099085, 126.9278056819142, 135.16395386601812, 151.63401132167422, 162.72556616674987, 166.34608622228234, 173.83491705059942, 181.72671801318242, 190.12708265468078, 198.55762353666833, 206.69428154106714, 219.10063953663786, 229.13736534689, 242.3177176748268, 247.69145846940202, 252.3368335028438, 260.0545730308504, 254.59464426881644, 240.97317883018763, 240.39451793331835, 240.6226149825478, 239.8768145967568, 240.10102572985286, 240.0805144103901, NaN, NaN, 18.825574219935795, 17.790518533631165, 18.19232090692625, 19.14509383955418, 20.282613881843513, 21.78850614900054, 24.397893729062226, 24.540561048884268, 27.000684928971847, 30.2321589340062, 34.643595436829585, 36.883192667713054, 40.03935517114805, 42.90229558854029, 44.62363362628025, 47.15181487552205, 48.90708981973823, 50.92402841227454, 53.16355959794484, 54.73789591978568, 55.829858545505346, 57.80731113480723, 60.516108511588655, 63.56349226785126, 66.75474916256749, 69.27999472746751, 72.35605367413022, 73.63185849682723, 75.49753802176545, 76.76436440046754, 79.21744014557618, 81.70913265856869, 84.99063304638558, 88.66106400042271, 91.07734909132422, 95.36031558994219, 98.77432827716191, 100.86327519846337, 103.38002724377323, 106.41774248111365, 109.57660424871645, 110.75363570442236, 112.96283924398777, 121.04388685658962, 128.23244569055086, 130.44375228226, 135.89914376671183, 141.96762512811625, 152.29849386305443, 160.12704245606392, 165.3529213300164, 169.98361635178827, 167.57345590011823, 172.3126779239936, 190.21594017514948, 200.7735553773749, 215.04116458753015, 219.87155350275597, 228.28744211106454, 238.84774429775936, 248.73363594938007, 255.88859723981898, 257.6466242974712, 260.0117160483364, 260.65287259545204, 258.98416588157926, 253.54523693819996, 244.93196672618012, 239.49869548845095, 239.13990613531377, 239.38928241327633, 239.65518259713014, NaN, NaN, 25.131704940531066, 23.838339820078833, 23.724150551022255, 24.788503813618185, 25.66978402195405, 25.224380008844523, 25.696274902681694, 26.685616039539315, 25.907977756215928, 28.405363651467475, 32.11636270108335, 34.170222300997246, 35.63214469190737, 37.39411084729208, 38.12154788114422, 39.954799478289985, 42.30168841819563, 44.57487871281549, 47.330081781942795, 51.00140608098293, 53.26936156374123, 57.30280538351917, 59.42517213304504, 60.375095680092016, 61.91180080016428, 63.00327225664808, 65.0595379600894, 67.99058285192267, 68.43096754506574, 67.17588075484726, 66.87573468461287, 73.02988974784085, 78.67974814498925, 76.9922127402339, 76.47619359502453, 79.85192238088221, 83.00881452723699, 88.73299989162004, 94.59473746866405, 93.34616581824046, 93.44036212527804, 92.15152987969475, 95.83681288988662, 98.96935771700997, 98.98128728687742, 106.3321519831939, 108.37843465749944, 119.6081927384241, 127.16132062160085, 130.83354148793578, 138.78446584683456, 150.5974522219493, 166.33344537152794, 185.79915555203445, 199.72739450536253, 209.43703040498397, 218.56202252694027, 232.84672780685352, 241.52924876242278, 251.53990362329657, 255.79704551181547, 262.95758600515893, 266.60827278274485, 265.56358857466245, 263.8599828166855, 259.7211842926021, 252.23524328887598, 246.78092503302832, 243.10052359431754, 242.7883108337979, NaN, NaN, 22.964113495516045, 21.634586385770277, 22.663230307876496, 23.94991763605833, 24.424181671438646, 26.629309194695114, 28.1731116956308, 30.157692006839746, 32.99058997652458, 34.53250931083955, 36.32950987514196, 36.28688272471947, 37.01991467235592, 38.634632735255735, 40.54354747536543, 41.863461376178215, 43.14607006097443, 46.19392597273978, 48.83584283708433, 48.12620093645237, 49.03893245733795, 49.83392857883355, 51.59473253999493, 53.21543597479145, 53.72761297477829, 54.08919976859391, 56.51070559423168, 62.81821588684363, 63.84351869602582, 63.09905876403742, 64.33517429899393, 64.54724250965025, 66.01086516969247, 68.35388842241305, 71.21233795464987, 75.98275840396616, 80.31532296345115, 84.06429978247529, 86.0412972638145, 87.20769464805238, 92.77698428712382, 94.54058599765641, 95.86449826755033, 98.67624375277757, 101.01873662860527, 112.33066498257307, 116.30734561596647, 115.13788801456143, 119.98716457155585, 119.57722816436069, 122.5301312747019, 130.65895952593556, 141.43903286453565, 152.6888427608502, 167.45927014011994, 176.6160504369605, 189.7451955513296, 200.03223589941632, 209.77244328976658, 218.29273147672856, 227.58554982914606, 236.01602991520733, 246.0216988752158, 253.01586284132043, 260.10850511093037, 265.52600677957656, 267.82177900468594, 265.54258464048416, 266.0786812941127, 264.64986524864634, 261.8962807388963, 256.1109088801178, 251.32482215682492, 250.74770346516468, NaN, NaN, 26.76348994453657, 25.727318610638843, 25.721828173243335, 27.00774734436872, 29.211961266821813, 30.567910041550032, 31.850708496281204, 31.771111119201294, 32.20872250617882, 33.19515125195246, 34.77015222769788, 37.080594475228196, 38.98380689274244, 39.52672360284627, 41.54114023438517, 44.58470759191572, 49.10485688138693, 52.807782650019725, 55.51126408077206, 57.155277601072825, 58.90362093888284, 60.29192719285828, 61.16331446647522, 63.80415304292154, 69.74098583064406, 70.6888279821524, 67.52862324412122, 65.77139262107242, 67.23224258248227, 72.8049126978418, 76.47201630460447, 81.38151695598151, 83.36346042370333, 91.44989523600542, 96.58460800794542, 100.53826415141425, 104.7912879654442, 105.97312174215695, 106.62792437494164, 110.08163956491853, 112.11188262866779, 115.21437022505923, 115.79273618169776, 118.89362465940377, 117.57476330308427, 121.68989993646204, 129.50421188454084, 143.069033582007, 157.71118812882642, 169.0232708591867, 181.23925566746112, 199.17718509121443, 214.20106030408564, 226.54112073203302, 235.60993268015073, 243.66925031333216, 250.79878061029476, 256.6658786802304, 266.100603394386, 266.0324684049069, 266.21924214443567, 266.12799035782047, 263.93499429088797, 261.28625343975716, 257.61062346617854, 254.93077926936652, NaN, NaN, 27.69308722876721, 27.321701296436142, 27.796417959299596, 28.010786806771353, 28.557633920192153, 29.54522561799966, 30.498858465282858, 31.340660569212318, 32.17748544834807, 33.27722279999499, 34.52393427906387, 34.77341681277935, 35.46868566028885, 35.866456944708325, 36.818526046740594, 37.617270718760324, 39.262821603425486, 41.795358324929666, 43.59128647158446, 43.4025516843385, 46.816279124782454, 50.488861499789806, 51.6574048639653, 53.116872579426214, 54.650016235345554, 58.17201239407545, 65.22022061268095, 73.36508822274705, 76.88167250649539, 77.75904592639571, 82.89655828627275, 85.97905219155285, 89.13157278784043, 89.49732550372146, 88.68378181823573, 87.86573862343214, 93.14108712304792, 92.99565698720079, 94.01028976772089, 96.87113560137433, 100.99434233141339, 103.92871834750565, 107.78446522354645, 107.59589767542326, 108.52382323374408, 105.77333323643094, 104.12895835152409, 105.79800311103969, 113.53180382609824, 121.08217220944489, 134.8581049628966, 144.45648184686442, 156.6721339338321, 175.51950029254903, 187.7986299949783, 203.68100610762102, 218.74501163276182, 233.04996401123842, 240.17422838061572, 246.23668940566722, 253.20360826286745, 261.41127614660996, 267.78671900819114, 264.7709963907911, 262.20754933161373, 261.28176216442597, 259.570046965802, 254.27801514631898, 249.61323854490044, 246.88693998538568, NaN, NaN, 29.827455128644413, 29.454558985695822, 29.74389401345914, 30.2520637239548, 30.982098938957602, 31.93365018702477, 33.403610043797414, 34.426303849406736, 35.48711520076702, 36.87792717500375, 38.37880378053908, 39.77036470625789, 40.829228204863405, 42.074391292276566, 43.31972121652915, 44.56578067060488, 45.62365018540188, 47.12217660031954, 47.26262020594502, 47.809943892034305, 48.3904912530729, 49.928783061684896, 51.765295746975156, 53.925120663334006, 56.304216913655225, 58.20708215396519, 60.30359261610947, 61.037681452449235, 63.0884808688562, 66.7606644377646, 68.99321006239744, 69.24550758282417, 71.84712223620392, 74.56416084116137, 73.93635383931166, 75.79898745970034, 77.12836885549859, 78.92883516170437, 83.48673531632798, 84.43937254880123, 84.9161355532648, 86.09752516683949, 85.80501215723089, 87.86153485516004, 87.12654893740633, 83.59619732623904, 82.40909744869774, 83.4308864986257, 85.62659409904892, 87.53481703850314, 90.17741046366163, 92.66384873206626, 93.4005756543077, 94.5739887842509, 99.27323213996473, 106.92360838468717, 112.67151389348092, 125.81032249178213, 142.94080342052064, 154.01978214187827, 165.0359821753279, 179.1048128831086, 188.7227678706743, 194.68666095721, 207.21762394151452, 220.9802564540997, 226.34428382792294, 232.23205073813315, 239.08935293578912, 244.98679018731957, 253.62414728555223, 262.66095406198326, 271.2157604255417, 268.20836787196623, 261.32965092271945, 255.35474821810055, 253.89609932337447, 250.5025685128104, 248.32634687320464, 247.4565484934748, NaN, NaN, 32.09002147723528, 31.79114201055676, 32.52590344270565, 33.66308341347584, 35.05782013142144, 36.04405788887952, 36.92070676380549, 37.68437912846334, 38.448706323909974, 39.43435541951649, 40.75381095625557, 42.25519914566479, 43.979414978178006, 45.25514771050159, 46.7566623803761, 48.96048256932151, 51.419484895937345, 52.33285679073815, 54.06126493641936, 56.70882986982932, 58.09700168820376, 62.27465010678043, 67.2727473684954, 68.7316461089186, 68.51252774100831, 69.09734493483403, 69.38876993187817, 66.88038678050198, 67.45783679148582, 70.90764900763848, 78.47060081584614, 81.05294290683617, 78.78247321033112, 77.53325881851003, 76.93532404626038, 78.32122539530255, 79.26641827907287, 80.13439371625758, 81.81563490701595, 83.12919840672878, 85.6527291175222, 88.03598978723136, 89.67943938247987, 92.23850717543002, 94.42760506358971, 97.18652230257845, 103.07614509763036, 113.57767851741997, 123.70901420214845, 136.6248364385308, 152.3054781801024, 163.95019505144973, 183.8094011281687, 203.73336121626778, 215.17596191587631, 227.80944914224062, 240.1667194494353, 246.42274485281337, 247.04365117617655, 250.99553317768826, 265.1203615322292, 269.5486427361328, 257.4300038977514, 251.55470574794347, 249.17661405053826, 249.0407121449695, 247.8708495201849, NaN, NaN, 31.683392429188327, 31.347443551015285, 31.969393597180186, 32.69823186866394, 33.39011221503253, 33.97048544798978, 34.66100612930025, 35.42510375960818, 36.152835963468824, 37.175658636808016, 38.3090202457831, 39.516021954528505, 41.130667137281684, 43.111816837953064, 44.83326897290415, 46.59196455395993, 49.051064811438955, 51.76656043421727, 54.00058745598457, 56.45904409434231, 58.62482057435487, 59.5079467031923, 59.28790113637347, 60.61049734714558, 64.42199412341932, 65.2319680517248, 67.42497517157713, 67.86400601068829, 68.01416983772687, 71.54368073885168, 74.34324356496539, 72.28630417430776, 72.35167752538827, 73.8221462951993, 74.25747563477601, 76.01913082864766, 78.8836872689865, 84.24609203359223, 82.99563339671371, 83.4273967415388, 85.253460173305, 85.97387993274484, 87.61476872412081, 90.3712316913608, 92.76772277445262, 94.78746319763066, 98.27637857627079, 105.81487608002497, 115.57447517700233, 129.41550172121242, 142.32134510801689, 154.71284205502243, 173.6099672443893, 190.8576908893167, 204.29160937096665, 215.33521705719852, 224.77129403627757, 233.3820555964706, 242.48310414816578, 250.51432381651438, 257.54355266561925, 264.88540864468183, 274.5623378245004, 275.0770201129301, 257.6481454624237, 250.02699812373055, 249.6864036141998, 250.0931833767521, 250.0694516971574, 249.49344194481665, 249.10359267546377, NaN, NaN, 31.31497106272985, 30.941832175764592, 31.52721961552659, 32.1815113540639, 32.946509867851795, 33.63536206505905, 34.25062720199403, 35.086644273305154, 36.292229534487184, 37.79190840349752, 39.550585235273424, 41.232939257016184, 42.87816698240942, 44.81861814131099, 46.6465043310144, 48.47539540362197, 50.04294079562156, 51.9073026407083, 54.509983756708074, 57.69935857808647, 60.66893610757869, 62.93611763753828, 64.18027106365297, 64.2481901171757, 65.27817492231465, 67.48231534859926, 69.6856636875284, 69.45536327847782, 65.34616918604912, 67.11981304022575, 74.54069651825499, 76.74464815522965, 74.76525686730064, 74.17747357091697, 76.74074431153977, 78.06395162109665, 78.50630318219102, 80.85875600269694, 82.31928386318548, 83.4816493822829, 85.97143032773602, 87.43080304623334, 89.6233727019703, 92.56488813798097, 95.14178473516841, 99.1950518425506, 104.88689808169852, 112.98875018667114, 126.44133035358199, 149.00119590701138, 170.23318817442092, 190.10800629860265, 210.30954677743995, 222.92844671703622, 233.73858437439415, 238.8215942456326, 243.8921807484052, 255.33621788386995, 261.2093836690566, 265.8024614796466, 262.54134889001506, 248.58201127237754, 247.35170405815705, 248.06511793525982, 247.88260893068338, 247.17303933536087, 247.15290491358218, NaN, NaN, 30.31556174087382, 29.722518532564855, 30.56756564318249, 31.4446973098675, 32.58233275004621, 33.60627921577216, 34.55595258842796, 35.32039071661771, 36.49138668351489, 37.69891027188058, 39.49641446784758, 41.58944711352048, 43.7911312437416, 45.40130986184979, 46.97377479416805, 48.655966835671045, 50.411654391808426, 52.27540223863598, 54.88275790194432, 57.59423053071894, 58.753613495294225, 59.61928469612495, 61.37310136816033, 64.74890014675964, 68.0450483203491, 70.23473373810599, 73.7598471967512, 75.96841763463632, 76.99172878665878, 77.364538655341, 73.03751708033275, 69.59075388872056, 70.10707648642331, 72.31746787367626, 73.93527429358387, 74.00465407286954, 76.58068565695396, 81.51511949544762, 84.0876383015575, 85.18748107936595, 87.26997721601346, 89.28011858375955, 89.827321634716, 92.21677776990505, 92.3999024171428, 94.05522891155617, 102.34045370152903, 109.67814384541234, 112.96256116291742, 114.77547177083878, 122.71995508834924, 140.44490035910422, 150.39121925665697, 169.47257517913562, 183.11015507992363, 198.03952171220888, 211.87394146367498, 224.3143290764998, 234.69665480684063, 240.02331961581527, 244.17013117891744, 256.81341039785286, 263.78866844276047, 251.04708248531946, 248.23730414535297, 247.2554471453139, 245.8263518579726, 245.800822047414, 246.03869315288145, 246.29884987595224, NaN, NaN, 32.910008922834784, 32.27833568680218, 32.90027110242337, 34.44370899284209, 35.43011283270054, 36.60132057553497, 37.585508525715156, 39.19979632584583, 40.663932608495756, 43.16475010594799, 45.77248144368395, 47.971963394456296, 49.98531332429777, 51.777174930150636, 53.34626670863937, 55.21096577445153, 57.18536719369933, 59.603171643764476, 61.4260686957624, 62.25272360542857, 63.71152530382979, 65.97555849903092, 67.35437354740706, 69.02981408006956, 71.29174861118999, 75.10421077448133, 80.46225071964868, 83.99429695181863, 80.40127171626308, 77.24113824557304, 75.8701350518854, 73.68591705281598, 75.30820347651454, 76.2654146629525, 77.58961620011442, 79.93146638409364, 82.19637358122317, 83.28549437918714, 84.67703958955084, 87.2406196232687, 87.95771124422374, 88.49461964637531, 89.76766258928969, 91.59162353713414, 93.78340852345349, 97.6361691898264, 104.98450976201619, 113.44725257449743, 128.9317446944312, 142.948236148521, 157.1774268410845, 178.6666286028305, 198.37176797283797, 218.1026313980898, 234.53625692765286, 243.63788194642797, 247.12171852770877, 253.34308061892833, 265.02566366783924, 264.21654944877986, 246.7916976060655, 243.9165772364817, 244.17990140092138, 244.57699700213743, 244.83688699886721, NaN, NaN, 31.388444606774023, 30.64604864783854, 31.046329408026544, 32.44257928697277, 34.318007651751024, 36.154249411799746, 37.767521663041144, 39.41833302490893, 41.401539692105224, 43.198394015520975, 45.55070276007592, 47.715683663165684, 49.95386163030589, 52.117783790807, 53.35548454570277, 54.33485992889705, 55.46202880417194, 56.47850427134795, 58.86549920752095, 60.69050940469694, 62.29687242263562, 63.973614374498766, 65.57498982474965, 66.66139679672379, 68.55737120094737, 70.22867390134104, 72.12148302674878, 75.63791599752734, 81.88691477758167, 84.77027235107663, 80.54433414358333, 78.15905239835796, 77.20872981249245, 75.59300066076466, 76.76481885637973, 78.22182880554364, 79.45965087553884, 80.9921574557938, 82.52182289274901, 83.38767803109407, 84.47456567842417, 85.12245182523141, 86.43752157871091, 87.30988263517229, 88.62371187151605, 90.81419068475779, 93.00503639466717, 96.30125758082741, 102.71035592521787, 109.54923749615021, 121.92634232198147, 138.5229999164271, 157.16785029460158, 181.6413988250454, 199.9146080498324, 210.42466661463533, 223.80297840625494, 237.73110035252586, 247.79748478236974, 263.39872852026207, 267.63376232555214, 250.58958734893764, 244.89371022182192, 245.00782144520352, 244.95130147231802, 245.1162269634463, 245.3664201207841, 245.629311073959, NaN, NaN, 31.165726826835012, 30.127472447862615, 30.639046312061673, 31.36794907332996, 32.3937467725737, 33.6777166867089, 35.47867193128366, 37.20382933152928, 38.81845398617741, 41.245825298405606, 43.63468573468178, 45.837789147417396, 48.26331119790948, 49.83487257065503, 51.85220587632646, 53.49934842692196, 55.476707398349824, 56.456724714551825, 57.399800856136785, 59.41771773396418, 61.72525083642554, 63.108452067793024, 65.37666046808954, 66.092169645594, 68.51171950187965, 72.0304497190015, 74.66140369556703, 77.58820335885785, 82.36600812358118, 83.36610138148262, 77.39748597660378, 75.41998933221203, 75.27504267345444, 74.67543202270976, 75.03369411837859, 76.49424949619487, 78.63030867638564, 80.90472257352845, 82.51268181981351, 83.38095104624018, 84.28389187074151, 85.29835016360396, 85.7964647845166, 86.56304648394739, 85.77941321072458, 88.8529935054288, 89.09900573213515, 88.57321839680867, 90.10009041278784, 93.68660627893696, 98.81681352594542, 101.89916148893134, 104.45642097701483, 106.50295212751085, 115.79657495910524, 139.82542723131175, 170.4387365595193, 193.83045049211714, 212.98414646768427, 230.09821507418664, 241.05917582350034, 250.54444162180582, 262.83510071747804, 270.6890514906187, 270.9568433384986, 257.91676053576333, 247.93524021330137, 246.46349804791296, 244.27575075215842, 243.91501708244596, 244.0884415393821, 244.2730740840563, NaN, NaN, 31.055557630507835, 30.202456385934504, 30.714434627612746, 31.814673304653496, 33.32041067879863, 35.232593343898145, 36.844989628312554, 37.60786159985361, 39.22140125162537, 40.3892211763562, 41.92858751664428, 45.205075189899745, 48.217679605565536, 50.52909928381305, 52.54221141676462, 54.002597973671925, 55.5357760069679, 57.14289152187621, 58.861726248962064, 61.280480654254504, 62.43998218620632, 64.48781335442095, 66.23606270257339, 68.72523474772474, 70.98608181922854, 72.06866460468618, 74.92534596823758, 79.61817268826105, 82.8503836327882, 84.17579615582795, 81.3470998834181, 75.38640744393778, 74.88380565673353, 75.1044992782121, 75.980278863568, 77.21794773740885, 79.50903084225178, 82.0025543933607, 83.31612816711687, 84.40268474829308, 85.01103520947233, 85.87420591052633, 86.15893762352674, 85.26513094830894, 86.71859434984948, 87.8768522135614, 89.32632029604173, 89.3119563430859, 91.06134851029923, 98.68289251515185, 102.19071455420162, 104.82362084382383, 109.82836448818728, 127.83942034600415, 163.96088911412744, 193.08074375963375, 214.62418089579535, 232.14279440614604, 239.95378518389865, 248.56798010542718, 260.1810175465726, 267.38753581497315, 261.8861878167376, 249.39311979198945, 244.58422135796278, 243.46451528846126, 243.75340449767086, 244.041420280437, 244.23210814712255, NaN, NaN, 33.64594586289366, 32.24044577760941, 32.899344942269934, 34.14746136666166, 35.802947823914124, 37.157933689795065, 38.62549320035493, 40.31363598242659, 42.07498386794718, 43.02008585238358, 44.671499138852944, 46.763793885342636, 48.89125381871034, 51.316986683000906, 53.627062486837175, 55.30935540405026, 56.80605027145806, 58.48767454466596, 60.093887798973874, 61.32817946500989, 62.491327510514495, 65.72082193784136, 67.02367145931584, 68.32937325907345, 70.30025481122219, 73.08191725706718, 78.07583233195511, 81.82642498112675, 80.81287035596736, 80.16082259355316, 77.76321738058729, 75.12585089100098, 74.68255751771396, 75.34180415480185, 76.14539822544161, 76.58051869632857, 77.98533792530888, 79.67635499435191, 80.6189314280156, 82.07674950511115, 83.27596218271424, 84.43843641217671, 85.30753785572746, 85.59030056346128, 85.58028725312109, 85.85637242321437, 89.07080957543725, 88.7592135102645, 89.33104602599846, 92.55116635332568, 97.83597462299271, 102.23121300183179, 103.97358107191478, 106.01869878381336, 113.67749285033987, 140.57570114849455, 174.93337357949184, 196.0145911066971, 215.18661803212268, 231.8575963715913, 244.31815687570491, 255.5055769689811, 262.4369324140268, 265.82204942086054, 248.45508096927892, 243.0642997304313, 243.5777700139025, 244.0879678442, 244.43537491770888, NaN, NaN, 45.15980647727301, 34.080872460515955, 33.0787629889868, 33.844594685675865, 35.38620102571013, 36.260713208373495, 37.134228192532234, 38.121082380121926, 40.328114782814716, 42.97648701096595, 45.068803162851545, 46.494965584002685, 48.144196267853395, 50.34621745472326, 51.99183626274744, 54.08345309228603, 56.06139518208326, 57.927904720792235, 59.90403897565767, 61.437303312861424, 62.748317071870055, 65.05558127690125, 67.13674465006093, 69.29285644938312, 72.11097686101967, 75.18792987296752, 79.73675105727237, 82.68521791402335, 81.77281410713148, 78.4394057190174, 77.31386087864668, 76.43722065256722, 75.66824789310398, 75.82440604744359, 76.0413487122382, 77.55217126075397, 79.90050103843059, 81.28987166304927, 82.89808012120282, 84.13178923847832, 85.14337406658527, 85.79409806260752, 86.6585039019304, 87.96232056911062, 88.60807505093618, 88.59072516845339, 89.90434949230372, 91.88054669775947, 94.07692290853046, 97.38282439500998, 104.01138466486113, 110.18730445232579, 117.03020105480103, 131.41642941721753, 155.39890966086875, 180.57636161543803, 200.69312637770355, 220.32393918610214, 231.82880330533874, 240.7786583691914, 247.23979583534796, 256.07979878678105, 259.4982707401744, 267.5696239944786, 272.29591771214893, 265.50444918451547, 252.4400833625959, 247.15492259855642, 245.04346709562836, 244.92175466282558, 244.9971006350824, 245.18530339886354, NaN, NaN, 34.823029933665545, 31.64402807335673, 31.785431259694423, 32.848229103571704, 34.0949846586896, 35.37597206047416, 36.54587498901889, 37.78938153248042, 39.03200051574412, 40.20149345335639, 41.888220514124, 43.905891186763625, 45.73683466793086, 47.34580310592165, 48.77020359976682, 50.71323811072122, 53.022825280619195, 55.777408823157735, 58.67573505060181, 60.50084909936472, 62.84398565252563, 65.07172875912887, 66.67174309571917, 69.41531221217024, 73.1168334440458, 76.48395161803285, 79.64027225727115, 80.85403795162372, 78.3056190345604, 75.2250149840704, 74.23646898796136, 73.02647317009026, 76.0041958222451, 77.37235545079834, 77.46994814458596, 78.15720033534384, 81.01896310120361, 83.25285522527463, 84.23047107662386, 85.0558106840188, 85.8471160496729, 86.49491111753775, 88.25069327127656, 89.78387697036328, 91.98072498488943, 97.05335606284655, 103.22233179564049, 109.61711638356658, 121.5487797194495, 136.3889034216868, 161.92046531463353, 180.38556975526643, 204.13664560343665, 222.56093944542968, 231.6075732874091, 240.48039784158868, 247.0749171861981, 252.52642671719434, 260.17707770995617, 267.52549768980947, 266.5741233930188, 256.81618011913474, 252.75992300987926, 249.01370047440903, 248.45607600660702, 248.6488560275085, NaN, NaN, 51.91673017421926, 35.67121821244097, 33.74526499746066, 34.03153784474652, 34.75976482719067, 35.78434063178029, 37.40008212143278, 38.717094793935495, 40.03604175151854, 41.944593897944465, 43.55521174683102, 45.16849325218967, 47.223498756793134, 49.12766854070001, 51.0294319652065, 52.193721196478656, 53.95030716362958, 56.88962116973497, 59.37844235486433, 60.9825153605851, 63.73195615986454, 65.73625873986622, 67.93020150831974, 70.6716000511623, 74.09075116337861, 76.06990997166824, 77.69329046800765, 77.5466936850165, 73.91649173152746, 72.23191703412787, 72.7156572623685, 72.11999962315295, 73.21671586751698, 76.30560724581954, 77.43744492201851, 77.95227306845146, 79.15649275704854, 81.49883366812499, 82.3718930266646, 84.97169631803337, 86.39141463741687, 87.84942292211029, 90.04005428188965, 90.94209843575608, 91.48953214062183, 90.9322405104939, 94.97126180466384, 99.73992254302767, 106.1739054929728, 117.757228541104, 131.04445202812033, 146.7510013140898, 167.4589515334269, 184.54586923366142, 204.51683608509472, 218.54176569951528, 227.15748640787217, 236.12319271471645, 245.79807978568712, 251.32985456325977, 258.8218101676789, 266.86751099842974, 267.3241683588136, 263.63913985980633, 257.5592947661353, 252.08619066964883, 250.98568746472344, 251.09157766731855, NaN, NaN, 32.50329625064442, 32.24033204794143, 32.82527551995867, 33.59117110763454, 34.43105527659845, 35.45465203236205, 36.58802743563318, 37.68482070651241, 39.00123901778322, 40.133649090762894, 41.56071163804159, 43.02414227695593, 44.524326080032765, 46.17121034563424, 48.00279373850686, 49.86948263556187, 51.88462785084255, 54.59896327080189, 57.34925224840809, 60.46861464022525, 63.290813907061256, 66.07547925705535, 68.67324897569618, 70.79496241046401, 72.0751577663838, 72.36789285033153, 75.49510585769536, 75.5424102889436, 71.32955607000488, 73.75566944515388, 73.69700073181657, 74.65389413701503, 76.52194538925083, 77.4798572246344, 78.43775788981429, 80.74678235273211, 81.69498712513261, 83.0840886927445, 85.27493957981012, 85.92100067341111, 86.71456518728449, 87.98782388640367, 87.61170451226963, 88.33756743712411, 88.14446978168583, 89.05345905167843, 94.74126315935219, 102.45334394344204, 108.14789490534874, 116.61821868212941, 130.0944831120008, 147.08884429637018, 167.80125725265574, 185.44531150605118, 208.64306259790442, 222.6742767897797, 229.04074068163806, 236.2693706495072, 244.25513054605588, 250.33863979065515, 255.44911420509186, 260.7929109601348, 264.0509445608782, 261.5444479832838, 257.7377013516262, 254.7031266934265, 251.21491957859638, 250.60914143285422, 251.01442761408413, NaN, NaN, 36.01215428696288, 33.53452485923902, 33.601529449940706, 34.405038421670824, 34.87560965154473, 35.78944456779221, 36.591244936157516, 37.46698536880114, 38.2687760058943, 39.40188776594399, 40.57133286126466, 41.92589734956759, 43.427255262804934, 44.92751356066545, 46.35320925844171, 48.29600118802958, 50.5325828683771, 52.73085784565606, 55.33422058528008, 57.899413705068156, 60.836055718829854, 64.02848539623629, 66.85013955452219, 69.08522716313261, 69.88432970420531, 71.57454148131919, 72.45445175081491, 73.15112147479427, 72.42164103087808, 70.70794520802306, 71.70817495727586, 72.437354704102, 72.20995150093607, 72.76131167471725, 74.5271503163428, 76.58587635592468, 76.84601033520516, 78.15790721640485, 79.43472873973072, 80.56895950799893, 81.58900650949039, 83.78580640854834, 86.3462537132745, 86.33275553241828, 86.68341147502379, 86.85032099485177, 88.12728552423565, 90.69632319852126, 94.17975875043875, 98.76953401648942, 105.75394793587024, 113.67237939345036, 125.09512958893275, 145.79471696414524, 166.28403143805988, 179.96495445399614, 197.68974775306162, 216.80314391434817, 229.57675776162927, 240.07641963943018, 248.964840118762, 256.74411959699796, 262.0687165021344, 268.21047086443417, 265.672171377732, 258.591468692651, 252.65840281017708, 250.5005005561584, 250.17975657408272, NaN, NaN, 38.52425767007105, 34.754071046445155, 34.78434386587644, 35.587439245432854, 36.86817861869674, 37.741223856965604, 38.31801991369174, 39.56175971628323, 40.98867507360439, 42.45204917696383, 44.247010823546056, 45.96671691230397, 48.05491055502414, 50.14229286164541, 52.34026682960074, 54.35131448245696, 56.65810164943346, 59.33420868117409, 63.30477952981197, 65.9779105156523, 67.5126992984674, 68.8642530009826, 68.09050978821138, 68.04809583622122, 68.12102076328704, 66.13256924107944, 65.50801146097206, 67.52384081592413, 69.208309412895, 72.14993391151688, 72.40906169431895, 72.6653550917999, 72.88665041718045, 74.02533889434102, 75.82479322235575, 78.10240007906125, 79.8995591815051, 78.90256401682848, 79.96029544212969, 81.27399300238211, 84.06338781958013, 85.60023100901812, 86.68893384322307, 87.78004525527848, 88.86770805782278, 91.51166493220074, 96.58033630307044, 99.44268812544325, 104.30042055794954, 113.35719352387046, 128.86342236954496, 146.56405922690112, 161.40392384298096, 179.45447488425378, 203.6139564065132, 220.26569688881827, 229.25049380402353, 238.11940096531566, 246.17958004229294, 256.0091847713359, 265.0988408844332, 266.792095366725, 265.57266462033846, 262.13068482641194, 255.59685031043023, 252.8374876224222, 251.59970762002348, 251.85217434377435, NaN, NaN, 51.1317734690778, 35.18541565029005, 33.55568156807962, 33.84247547409337, 34.129276130928474, 35.15514818354177, 36.327709894272594, 37.49968337327512, 38.967744380796056, 39.98993210309952, 41.012837341209874, 42.183941478488855, 43.35353844244724, 44.966637715870085, 46.72599413566199, 48.33710907851832, 50.390939774571706, 52.59245877893337, 55.236444525534175, 57.58296987536917, 59.85701805803429, 61.76692489418739, 64.1612167679973, 66.73135781034082, 68.11988214067023, 69.18010794545731, 67.96608043870734, 66.0957618428516, 64.25203351298113, 64.44154227942073, 65.28420983075813, 66.59542958980929, 69.93517385429583, 72.94717834468014, 73.8592478092067, 73.04931248921379, 72.97312461129154, 74.66044670742902, 76.19502752343347, 77.58433347287874, 79.23271505808647, 81.43227286984636, 82.08579588967633, 83.83878393198502, 86.0345168913596, 86.90691987883751, 87.7720017536275, 89.5243265075933, 93.04528688528714, 94.79736032216337, 97.44741165377378, 102.7479710546618, 110.91870590457589, 121.52433980236779, 133.24665836757336, 150.76090816118753, 169.86137399279963, 193.31984318918705, 212.32832127159506, 222.9025578498131, 234.1681757983189, 244.8843161025506, 250.25082539185522, 256.72889732700895, 260.8674731944062, 264.84356468880134, 264.49444821915654, 256.8311509379599, 254.0435440703565, 252.0588437017123, 251.9915140436925, NaN, NaN, 34.262879074662706, 32.634840261705335, 32.99873413082677, 33.58152876554952, 34.0889171552317, 34.966026195543975, 36.28552680598321, 37.19781105228635, 38.18371496213357, 39.17033086902794, 40.52584366461859, 41.917966597706325, 43.9376031945736, 45.3640982003088, 47.12281237451112, 49.21401726615635, 51.413391201133976, 53.46605283867503, 55.22179343712757, 56.50193840938636, 56.49664742648443, 58.994225884809445, 58.62325988176222, 57.44468277398659, 59.72076670920724, 61.26629318224823, 62.58013724075413, 63.90752660543854, 64.1995393432148, 63.98007736353169, 65.66727976730911, 72.50411728460527, 75.22509731715753, 76.3347719291531, 75.22394807091786, 74.04248187676001, 76.0319000399295, 78.45567109430415, 79.84187177895353, 80.57012927256052, 80.78020867483043, 82.79503677098674, 84.06661966168299, 83.13785390871318, 85.14723791905192, 87.70447595799264, 90.26888084876519, 92.83272990898523, 94.47319159297162, 96.30702754480168, 100.16992227525475, 108.07475204072003, 119.13400007750474, 128.53154455213084, 145.72041548435033, 168.68605877896505, 190.0265902494059, 207.19671568300652, 219.5719738598131, 228.81614162940375, 239.20566281022124, 247.7521440634587, 253.73582960664862, 256.3872976917702, 259.8825285240161, 267.5555817359507, 268.4117130288364, 267.6813282519468, 267.0502406982261, 262.8818442091029, 252.41071017337492, 247.60378085678587, 247.77432352765913, 247.96890946569792, NaN, NaN, 34.33852377103652, 32.52595127501537, 32.77759717283, 33.98756866543055, 35.23217142497529, 35.77563145494105, 35.438327452757996, 36.02031863030415, 37.66941526169175, 39.54080144844602, 42.36842660265105, 43.356731543840226, 45.815646075966995, 48.20291313355413, 51.3693065459967, 53.34854572109285, 55.07535676734086, 56.79932296082183, 57.85328822551961, 58.91330949540136, 60.31622295714637, 61.707836523889775, 63.69137585857366, 64.63985820195988, 64.56143059208539, 65.8128972307363, 71.5469558838277, 73.59519983513275, 74.47188281362942, 75.71798528832359, 76.67709595476249, 75.78918527010337, 76.08351639334938, 78.3605779614949, 79.16604086818779, 80.18056251843268, 81.49481847464101, 82.06945316010267, 83.01407260439399, 86.38436207467096, 88.3527557466077, 90.5535369976915, 91.6437831270014, 93.64818097326888, 95.47809742595119, 101.17697718151335, 111.86532482888475, 127.17763364057251, 143.24344956778583, 159.13139660351658, 178.39297209458078, 197.9623654267403, 215.56536602544654, 227.387203688999, 233.79544470470145, 242.23330869889654, 246.40115473565092, 251.93204083691734, 260.94095283507534, 266.36108606180215, 267.4791169606709, 267.1619808264426, 265.27304300938545, 259.6228829714854, 252.33705688826925, 248.3926185703824, 248.3425618151838, 248.53574318892444, NaN, NaN, 36.739289887330884, 32.9711643945451, 33.40985692486786, 34.434979734917746, 35.68193903245394, 36.99995873515272, 38.058284333936854, 39.11841394599556, 40.32610313059294, 41.64688288898765, 42.78112569791842, 43.54492617942311, 44.752822202111616, 45.84871937705973, 47.28206652475435, 48.822590285754934, 51.06482465938983, 53.2641937036108, 55.539300426903786, 59.36152219202791, 61.34633298135983, 61.34039327130184, 63.027913017582215, 64.41138466844868, 66.0243686894151, 66.17020537424322, 68.01072312184597, 71.9157863829423, 75.5876302811044, 78.60382656041139, 78.82458241362912, 78.34028439173507, 76.5601151924476, 76.11492845466809, 76.8418336983604, 77.74542148123845, 79.31953961087825, 81.10896222342669, 83.37119994224072, 84.79560458761023, 86.87683368772846, 88.18833066868253, 91.04770579025211, 94.79228761157789, 96.32353811322079, 98.52013130841497, 106.47062711072624, 119.73475982367884, 133.9057856706273, 151.8599695235672, 169.3865365633006, 188.80254713959175, 214.43770015752406, 230.00382945233198, 240.88394144471803, 247.90819544071087, 254.8058696355194, 264.98866890360114, 266.87685425064564, 267.5025427066237, 267.57043272981224, 266.63910179730203, 262.2227376989662, 252.25050907538468, 248.36370026964892, 248.41612200464135, 248.71760783912006, NaN, NaN, 36.67058592712896, 30.169717571149484, 29.648865142845803, 30.968878781863776, 32.069258354898146, 33.53629625952673, 34.92713055006752, 36.612211610242106, 38.59326325136166, 39.46818147135966, 39.89979391309554, 41.586040677404, 43.64010358761106, 45.693374039067905, 46.933898593169204, 47.81330192641036, 48.689032329992564, 50.741438789378606, 53.16348735319967, 55.8812145808991, 58.11840436109902, 60.319303500879975, 61.93006220532172, 63.20916386464081, 66.13980308270045, 67.27892014038937, 68.27122224203072, 69.99175532015909, 70.83557188251947, 74.1063725665554, 73.62898242733154, 74.94982977517107, 77.59625729546241, 80.02538409431556, 80.68207157849739, 81.6651572301745, 80.96907317829319, 78.64863605267008, 80.1146509728737, 81.10416867826795, 82.82058338929883, 86.1947927512526, 86.92650116142387, 89.70856358031999, 92.93433392731914, 95.58451646517922, 98.08646237106278, 102.93629024067404, 111.63075908914209, 124.30662084862372, 138.03279991959855, 153.97909584353914, 168.76160065093396, 185.83046619985052, 201.2135228879662, 217.5728527448446, 232.84951242396914, 246.35897163420643, 252.8439966358014, 261.4231965811717, 265.8974765050644, 268.3772724173144, 267.4707964970133, 267.0891619457841, 264.91776450215946, 252.68187442565204, 247.94969671057711, 247.8031019406022, 248.20577718613006, NaN, NaN, 30.348742405552713, 28.16867061047757, 28.49511376358156, 29.41180575780752, 30.365681443946716, 31.31952728958485, 32.86063206668966, 33.85178414247405, 34.875734304257044, 36.74749241580549, 37.36529393585783, 37.945985217791545, 38.67624262879984, 40.14238102959593, 43.29825312723023, 46.162162930233876, 47.739649169555406, 48.87123320221508, 50.96229831297883, 52.320435267014176, 52.610056033324284, 53.379333952724394, 56.31073855882548, 59.61357967347791, 62.805329021021905, 66.47959358720176, 69.63147530002296, 72.82867848491034, 75.64417934323407, 76.44422108022933, 77.43102132790602, 80.1101297921342, 80.31833943876487, 80.83297141553861, 79.62737863621015, 80.91274652094741, 81.93478996634131, 80.76044940362307, 81.04675628358235, 80.276844354499, 79.61818567460695, 80.64291413112882, 82.6910756512115, 83.41864862290159, 83.7048732097865, 86.33720247964978, 88.97666491753913, 90.29499935803376, 93.23136715783842, 93.81272199088745, 97.33093924396762, 107.33120827089164, 115.86714316525664, 127.37882272954785, 144.50320929381996, 158.54080249311207, 176.01869989668086, 191.48337576353893, 204.11240197729623, 215.0879752390339, 225.8624805217543, 237.95987954675405, 247.80597139334282, 256.41148197158606, 261.8248168315665, 266.09435142799236, 266.9101197663576, 266.4441134221939, 261.75057584741637, 254.06707062847192, 249.89647052752372, 247.95026927207988, NaN, NaN, 29.950680886926456, 28.656483008397075, 29.316028281744465, 31.117844054769694, 32.25499349223071, 33.611713890642065, 34.450182464281056, 35.144497934129305, 35.72870855795814, 36.313307617928245, 36.491474972578956, 37.84533757902916, 39.68107531279759, 41.585750678828575, 44.48779623491082, 47.27813938644725, 48.85165916019006, 49.68845587101894, 49.86696112633735, 52.58361219501801, 58.05942311839072, 64.44839132735899, 65.17974331943888, 66.05227755306977, 68.7660772080461, 71.92845427020177, 73.98861639879776, 78.61924720596129, 81.2593018273514, 83.16985232115803, 85.43675611537032, 85.36394286766183, 83.30166737749391, 81.97284863869706, 81.67525314283674, 82.7796482954842, 83.65542801118195, 85.11504690311594, 89.37655027122246, 89.8087222893382, 90.82842224934012, 92.43413387311165, 93.45482967417193, 100.65240706030663, 107.58442006677815, 116.13961707088313, 133.87812337851727, 147.0114019696071, 160.16607400386235, 174.38183016003666, 190.72418902875572, 204.11762794484207, 215.82449389135562, 230.57534540432545, 236.76971604938484, 246.17108952343614, 253.74294064928796, 259.3507183593953, 262.9493737691629, 264.63184397158983, 265.33353884758566, 264.0817823979605, 259.13684589882183, 257.1473870935725, 253.17749489218863, 248.54533222348886, 248.13997785617204, NaN, NaN, 32.89493370169752, 30.567843587599715, 29.64292213467525, 30.338383412801637, 31.65893578892389, 32.870202289030885, 34.006941640233535, 35.03293423658797, 36.42574133354608, 37.194863647011566, 37.88613271921641, 38.98456837550121, 40.48536021235354, 42.872481146437664, 45.92235312775038, 47.64249282048605, 48.22100714391904, 49.42527285209523, 50.44689166694869, 52.0571591210003, 53.92649517340292, 56.20125776304252, 58.175439251383935, 61.18169709033727, 63.22707049134655, 65.57110670021642, 67.69598693628129, 68.79337550968995, 70.47580071653341, 72.75086586531654, 75.25152441745118, 80.4662190891116, 82.51556066999918, 85.45780441040893, 87.00054672212906, 86.41513418402488, 89.7164576265294, 92.42544853195982, 93.89107202659078, 93.23611803502268, 93.63828372760025, 96.3927655871533, 94.18685383099955, 100.2409304254491, 100.79991607822963, 105.57018674478344, 115.49873087616729, 123.97412887954133, 137.2856613050069, 159.49971862897212, 178.7731251364426, 198.16682811986087, 214.04837059219776, 224.8919945886474, 233.38139144348062, 243.64404597652688, 251.70981430774296, 256.6575639178689, 259.0495477615819, 260.0723247187183, 264.5428928118693, 266.5111122339867, 264.5443452737095, 259.12531423721254, 251.61564935286373, 250.33244513474955, 249.01783831480768, 248.845203055696, NaN, NaN, 34.77472301319023, 30.272019882596922, 29.901824250395574, 30.634915173086036, 32.547929593951174, 33.86597675229869, 34.8923072139076, 36.91553137378167, 37.71733126413065, 38.41086428040415, 39.58515131020383, 40.6853562989706, 43.365391022895984, 46.07998506055057, 48.684643692528944, 51.66189543078722, 55.18770416394941, 56.17232075180884, 57.05156122687263, 59.98836662819903, 63.44491136165922, 65.42012562513716, 66.8880372031426, 69.97132553302069, 71.2838707649608, 72.16499845108068, 73.99744854177084, 76.27092441411234, 77.58919034412857, 82.06252673043807, 84.3465019557922, 91.41116642133166, 94.49645248159601, 93.75881811213745, 95.81236149492942, 99.47393368311516, 102.55439863830814, 102.62387699756373, 102.47727365186824, 104.02325442469089, 104.12986926383657, 105.04883199491877, 106.69672596256804, 109.45727945772269, 114.41918907426218, 121.4063396492537, 128.77986792187352, 138.36520243758994, 155.04704806639106, 173.94265212054557, 189.33021208583747, 201.80069923827807, 210.56454824388436, 225.0682733461202, 240.5928914916674, 248.2921450922541, 251.95613069968184, 256.8081452145644, 260.69043489675664, 265.2796866647047, 267.3972280906039, 264.76071261044336, 256.30089739432566, 252.2280645121218, 250.84638847943867, 250.30760935010892, 249.82260472708722, NaN, NaN, 28.204419183048643, 28.27598739182182, 29.452734777326796, 31.291426420886726, 33.42515454582815, 35.48244526873472, 36.359024527925655, 37.08803354497802, 37.078110450568225, 36.85392430739635, 37.06920768686347, 38.39004195597616, 39.70981578998093, 40.733208462944056, 42.71373992186032, 44.32734082655062, 46.89720010211287, 52.484954512403235, 54.984572227614855, 59.4632407734596, 62.62376837866473, 66.15502321405455, 69.01499642061654, 70.99879867067135, 73.63408255457765, 73.25962530330015, 73.09803885884035, 73.82877599227184, 76.31361336965891, 77.70743625595838, 80.64146613308428, 82.76130254302167, 82.90185733777048, 89.14319100031024, 92.90198517696105, 90.10195247116279, 94.65985607879992, 98.99868680062077, 98.20063330769773, 100.02627155910547, 101.63864156059194, 102.18872341276479, 103.0919266723618, 106.21635952008303, 108.80314595124834, 113.22273997018715, 126.09235067820593, 134.9549844685848, 141.789497290711, 151.9598095025097, 167.909452306315, 187.79870428611068, 203.26988173232942, 220.0754496495025, 229.21434970538294, 233.6666020586287, 239.4066085320926, 247.7496023793832, 251.9482659720034, 256.6146826836982, 261.6285182787181, 268.76622665442704, 266.4260954562535, 261.7767198014735, 256.68376944581814, 251.31702547929697, 250.342126741569, 250.45093546750147, 250.78110053297607, 250.67505793013902, NaN, NaN, 29.344310585554112, 27.348923916121375, 28.156192673462638, 29.47629482568458, 31.09293306755753, 33.37128490211201, 35.72087741673162, 38.00108530998992, 38.58632894686018, 38.063639426457314, 37.687158889042124, 38.49131312791784, 39.21784898438918, 40.23822156619713, 41.40799515940624, 43.093847192056764, 43.97303060987014, 45.51126359277563, 48.665532206582455, 54.175412759485056, 53.54396997870787, 55.223466258433376, 56.98174541030652, 59.54943015962707, 63.94973825594138, 70.71012205985727, 74.37927338970194, 77.59745603342387, 80.75369584686615, 84.13470870027963, 87.51384431081064, 88.24129784322727, 90.36710238484243, 91.60834526587651, 89.90893736186443, 92.40121924915897, 100.11251862270458, 105.91516879621304, 106.21619206199863, 105.61653497213864, 101.82067779744422, 101.45855737620266, 106.42641902535215, 109.56670116599436, 111.2337370242519, 116.02179478675966, 125.06574387263079, 131.87856913959092, 140.58322008824965, 160.03383034683026, 177.58868438272032, 192.68294151308825, 208.32151893018505, 218.05207680641118, 229.71284929633458, 240.2141762784856, 244.83598963906215, 248.11122686456437, 254.13341249246167, 261.32799961214636, 257.77157181103297, 260.88250375093304, 262.0197502930601, 260.8803904524508, 254.71780255927516, 250.70726448798084, 250.08647422396388, 250.4087831205672, NaN, NaN, 30.91089524319357, 29.39467423582652, 30.829210910548763, 32.22554592400043, 33.4022059748084, 35.38663550722963, 36.930597166194126, 38.39731446553491, 39.12730603507649, 39.967050087414975, 40.80644483992301, 42.12532723688825, 44.14030675058558, 46.34243818215392, 49.424333648155084, 50.33705640216491, 52.5756555244249, 53.41630390527763, 54.14861638051368, 55.20760509154346, 57.11570912096584, 57.842750198341776, 62.321588203517884, 68.55601090018031, 67.95690467574033, 70.88901894096533, 75.80862391362787, 80.58149609300023, 83.88552270753833, 86.89276154316897, 87.70435313276342, 90.19582271418588, 90.41801536836293, 90.05020854509316, 93.1315526575578, 97.23090710114406, 101.34283707570648, 104.94434697015551, 109.42549360941622, 112.50262146393328, 111.37529739266108, 115.79530164611721, 112.14627366351212, 119.15077774809066, 127.64478544851961, 136.32416793021227, 144.6212020810981, 165.7283989422765, 180.7315112245882, 191.85685382354933, 201.62585088984827, 221.41623861003336, 233.09322834513597, 239.58284814622476, 246.18312867700652, 253.38916397011442, 258.6589197371901, 261.45806823653237, 261.9314283919187, 264.62431481495884, 266.2599919530258, 267.2490140753673, 258.3041926817653, 251.26626387476253, 250.58946243806267, 251.10078631093364, 251.39407686286853, NaN, NaN, 29.3906830017219, 28.280025765599678, 28.49729242458693, 28.714217343946363, 30.1105920949601, 31.615961831044498, 33.04846552738428, 33.89249483890869, 34.847237832026615, 36.94472149860481, 38.77943267006252, 40.39168548557354, 41.01097266915071, 41.924040855272075, 42.79863609496476, 44.89231124853754, 45.94646257785686, 47.85409241641305, 48.58080229282667, 48.099473863307345, 52.688479142949156, 59.23199426555484, 59.88647341429239, 59.14360786496564, 58.767387390995616, 59.78848276187809, 59.710534736519755, 64.9227723137807, 67.3467604404159, 70.5740254934724, 76.88578783318684, 81.51063293951152, 84.79973904929712, 85.73663916969367, 89.99338744653966, 90.50810557172152, 90.72745325962966, 90.21327127273852, 93.52253274595404, 94.39421230401078, 98.11066324532074, 104.37583339288153, 110.0695994103557, 112.99788239808407, 111.35972247414584, 109.71802204807186, 116.18161653494305, 124.13582721187028, 135.95573953308718, 142.21428092988157, 153.70808809547157, 173.65641403056708, 180.9146016542522, 193.33129160201526, 214.42266319948504, 229.7381563564433, 234.654874126723, 236.75755905625957, 243.67926407754194, 254.97375937300134, 255.8098796542776, 259.67219942647233, 261.8867351499456, 263.1155846831427, 264.81379423731215, 266.2598617862924, 267.67596786368244, 262.50289995939346, 254.21874940899406, 252.16407318639202, 252.0682268892406, 252.39565580978652, NaN, NaN, 27.065057154124446, 26.764161716415213, 27.53481026537697, 27.603354024626167, 28.186082188886616, 29.69376534786583, 31.456169413742497, 33.182279157244835, 34.94562851171694, 36.488794800676594, 38.14329686985148, 40.421461287234926, 41.48260204881406, 41.880820321116644, 42.72006006738944, 43.85404977921425, 45.249617674872844, 48.517992668665435, 51.967705724700004, 54.4992756789453, 55.85122061427953, 57.535328912538574, 58.93155210616161, 61.20858931044499, 66.93933170755841, 73.63180105893746, 78.76584797262876, 80.95996172535332, 82.79189968305184, 85.27613877185833, 90.33367766361295, 94.80245240693039, 93.4117062233599, 92.02269916365785, 90.98400954163878, 92.29703931631684, 95.68428224207055, 102.30677100938308, 105.08167265397293, 104.34020350033039, 108.91526303432745, 111.56580067687672, 111.80904192540898, 121.13290675423495, 131.77239578506888, 141.0903488595326, 149.7001980579794, 168.7773963412649, 182.60356472830745, 195.5148099059472, 219.67671722138306, 229.54342373106448, 235.8968110019359, 249.7491088981033, 256.65678829121947, 259.78642447876166, 260.77335521300233, 260.8119620812434, 261.594666040069, 264.37179382163794, 266.3952337993557, 268.40573285411796, 267.0226877180711, 257.96759876814787, 254.9543642869718, 254.92369969984446, 254.99616382555627, 255.1723251547375, 255.37685082345575, NaN, NaN, 25.3746197408656, 24.337985360511706, 24.88613171592938, 26.0234369248167, 27.602985722048494, 28.44393634046211, 30.613471202091265, 33.00411097742049, 35.69055795100971, 37.56324827780582, 38.6990719509699, 40.05685656418298, 40.74982011318011, 41.66274354805312, 42.168270262087404, 43.00567191263895, 44.32367573776685, 45.34920072204572, 46.260518339014205, 47.87006531216568, 51.46876816375695, 53.89188109124194, 55.209255219537184, 57.51637230675087, 61.373351474109036, 62.68440576245977, 64.32656637260457, 67.18427322241173, 71.03497468876881, 75.9998160599481, 80.40474856817941, 82.3805544624006, 85.13566299924584, 88.55703422561756, 98.58472888931105, 99.46681508652003, 96.26557865894937, 107.83991640789716, 112.92827642152552, 113.3821697826291, 111.9281824658814, 111.95041548865085, 120.39433004851124, 137.5350095641768, 148.47004473515938, 156.46169729929483, 166.45793158076546, 172.39471056572995, 178.28410854259675, 197.5029919195193, 220.14843416811877, 231.05747817297376, 244.59000787112905, 256.67914451718536, 259.07645505372443, 260.0551232097085, 260.69406010685765, 261.7434305625877, 264.1195236081656, 264.14709042244874, 260.4163140595703, 255.97299690192594, 252.4582354809795, 252.40712552575002, 252.72833831894914, 252.97818727770326, 253.0756772961405, 252.97192652561867, NaN, NaN, 28.02142162214453, 25.991229061872893, 27.60648273812048, 27.89546536687357, 27.484290479867813, 28.61835739777716, 30.306608237205044, 34.05885035173562, 37.95603912878472, 40.4520605725567, 40.9598985309769, 42.13306981962367, 45.43704370846285, 47.82406628495125, 45.46581057664579, 44.941387916401794, 46.40593585159415, 47.97876282053871, 48.815968739556205, 48.953695498363885, 50.932457485813885, 54.35278744752852, 56.56143061717877, 59.749951787009, 62.82712257244782, 64.46804950532055, 66.55131200142834, 69.85173504547573, 73.48260740259953, 79.75944978606914, 81.51907960838646, 83.940532659968, 87.24774458612369, 89.78231179850103, 97.59356701193651, 104.65373386244303, 117.10408470263928, 117.77936525480021, 113.92026321926046, 112.60915531326758, 110.58435796726967, 110.61557396432214, 116.81771954858566, 131.8394529907877, 143.17358273230022, 150.3566897654903, 162.2067962663, 175.80293540681532, 201.5187614902775, 213.40131337852347, 224.60617411555526, 231.74793477415872, 241.2675121301503, 245.14421214685657, 250.22463892675506, 257.9349207674198, 260.7384242465362, 263.3976798262921, 262.2876066410975, 262.18798465330224, 264.0262897780342, 264.5140541788742, 264.9556291948502, 260.5636027753833, 255.98286299461506, 251.19611675481218, 250.28068770645075, 250.6059703313501, 250.71804975182255, 250.9746080078453, 251.08881536934578, NaN, NaN, 26.76856750016089, 25.32877648974365, 25.80309366553421, 26.90357863395794, 29.955673304339175, 32.60614515004919, 33.70591759472315, 35.06421896555176, 36.273204673489225, 37.48367025040769, 39.765009020890304, 42.07794761153275, 44.94014680337327, 47.843322590721066, 51.480115348012006, 52.90732072198371, 54.29195921243125, 54.50302963106752, 54.720088671912265, 53.72377946646015, 55.59283255251073, 56.134239119671186, 59.21035051682415, 59.75475684278233, 59.302735414161056, 63.925713570626336, 68.98811504352943, 70.4132547665286, 71.94676223977565, 80.86127902539634, 85.92368543586042, 87.0381766295346, 93.54463243552011, 103.12053483781668, 103.45526094726924, 101.90548165514365, 102.90375763604625, 103.69537911732408, 105.13775476409144, 111.19772451872194, 116.69832198670993, 122.4558401811945, 130.8477796499813, 138.60906700523208, 141.06887235280945, 139.30602342447065, 152.91177509020892, 177.88224201762176, 206.06277286846756, 220.3386216263845, 226.86255170427182, 231.51726522146484, 238.74137101036985, 245.1702987267106, 251.59923085717526, 260.5906692459555, 262.8232644911844, 263.99487283218326, 264.7135661460247, 264.1145198261076, 263.3405739567716, 259.91054490280555, 257.29026308107194, 251.6050525532619, 248.23752266021106, 248.26364541432352, 248.5177914604486, 248.76702837247973, NaN, NaN, 25.775838582447797, 25.73558943323872, 26.544582152314067, 27.867550257837856, 28.821212286585563, 30.141300487549717, 31.277027296368615, 32.37657618264209, 34.13881202165719, 36.6015378527773, 38.582402321290765, 40.48675157979866, 43.166841029201116, 46.07136965091851, 48.42033290579584, 49.809693739971735, 51.78618388399232, 54.46668153867915, 56.33843046616094, 58.28454198551016, 63.788949522649546, 64.22344054790823, 65.65164805604516, 67.95552289366488, 69.59622543316587, 71.4569380735104, 75.42576228733073, 79.06025436385809, 82.46674737681798, 87.08991377481284, 88.2949907144124, 89.17092138171547, 88.50498535127096, 89.71039492194663, 93.78892417539534, 96.44032455070942, 96.90233056724603, 101.77420808370559, 111.91150569022629, 115.01434055834652, 123.77464342959125, 131.52156460144028, 138.24538279979348, 143.93953277711233, 141.35148993152384, 149.69906015059135, 167.68962637548705, 195.7720918208695, 213.52619151059122, 225.9049738467965, 234.97905331167965, 239.0085740329833, 244.77832576454898, 251.48964225500842, 260.6855886772097, 261.48686563619316, 263.1385954142184, 263.11062110534664, 263.9749828599073, 258.28105917842475, 256.5890045224235, 255.94585518040765, 249.5097169180364, 247.98752533673365, 248.24322659502317, 248.2741685910718, 248.51761556154761, 248.53405637128583, NaN, NaN, 27.475356939913123, 26.843791135871673, 27.61304060131686, 28.381638448972293, 29.36994348792098, 31.13404794597969, 31.829234631244773, 33.554080741630344, 34.50892167123228, 36.6727489061427, 38.32374340121133, 40.451323082479725, 43.35037867934392, 44.268895598124786, 45.69461463755858, 45.86937178586535, 48.77210403803316, 53.075300336481504, 56.67501732398095, 59.46147913740105, 62.32212317286818, 65.1831134769405, 69.14657940417999, 71.89604858876686, 76.18678890063346, 79.1582766124879, 83.0105487464516, 85.20838714403187, 87.51616083018342, 88.05103465756704, 86.07341391986547, 88.49658343206346, 93.54793611227068, 91.44243804204599, 91.54743838385974, 93.41580515363205, 93.6335144978924, 92.19590069214057, 90.76959668674132, 102.23133799140284, 115.12312270970473, 122.8614273098745, 121.56268407778904, 126.89551041433704, 132.88064643811603, 137.76947185323127, 150.4105110443259, 161.07932032463037, 166.39112018647234, 169.55637112695095, 183.24143473334036, 209.4602151059541, 227.22909179557803, 235.4994249412514, 242.17860529362778, 252.4151515536774, 260.0275060830699, 262.002822840847, 261.9801843753621, 262.984762376922, 264.51763556077793, 265.79667235561345, 265.6353503783549, 262.5867971650239, 256.8529704491016, 254.93551060751534, 251.57033953195304, 248.11167287404527, 247.9991656515376, 248.17705815648546, 248.34892685984227, 248.43835960514843, 248.62468367976257, NaN, NaN, 25.47713216015721, 25.068868023933923, 25.72853848101566, 27.972932316784966, 29.738564604229186, 30.579119559636954, 31.60483925375729, 33.88429794797032, 35.090764636047744, 36.22764694108948, 37.83944540049761, 39.59827045498865, 41.57405176893084, 43.00257955046995, 45.279839384408646, 47.95840046221004, 50.30767036050717, 53.35632869407, 57.02882626835944, 59.601300222274354, 61.24662171854408, 63.14387861285935, 66.66400788987737, 68.11755825625013, 70.6085344580198, 74.42549694140696, 79.25918625288399, 79.54142613607077, 80.55720437002371, 86.57517661279088, 91.56738545428618, 92.15063633110316, 94.04850582787941, 91.26655729537323, 95.37342952131306, 109.31953309867498, 115.34033238798563, 120.9467100305031, 127.42423550291015, 137.06356736273298, 146.3081366637691, 155.34280683736532, 159.51303303223094, 157.83527229091618, 162.77834847070656, 177.6529038468996, 192.55300334217785, 201.70520996702996, 218.07029875112303, 235.04747732101407, 244.563205529786, 252.28490969191733, 261.25526188125093, 263.8416014151932, 264.25507055440477, 263.6459344875968, 265.7914295153785, 263.8762267436324, 256.4247499380388, 250.62732217189648, 248.0806772477884, 248.06803981279342, 248.28633962219186, 248.3889293689058, 248.52382083343971, 248.5815921911626, NaN, NaN, 27.4413371438828, 27.29085241702471, 27.508278002490496, 28.314516827106278, 29.96833618381884, 31.364974176463704, 33.35103469084179, 35.039621823508995, 37.869442464798816, 39.59230695837892, 41.16962664216967, 43.044560294895824, 44.88693069506303, 47.382443069412446, 51.90532214204061, 53.73828067290166, 56.011395717315416, 56.14995903148249, 56.65952359973792, 58.7874823047104, 62.71071648698952, 65.78783052834646, 68.53549114330218, 72.83145328054114, 75.0252363483373, 71.70635131264532, 68.17283623618872, 76.09621215031784, 81.49121545794027, 75.54630545673328, 76.97059366964, 81.03230587465927, 93.68684542412106, 102.71322501637309, 106.5735471267478, 110.32434940932197, 112.95832941449798, 114.93544973247604, 117.23678060001568, 121.98309221618445, 127.4179711339016, 135.98617692606166, 145.63209815463165, 153.78546375743292, 157.7802931297863, 168.16531366519462, 171.2561591815013, 173.64852086934056, 183.321984987941, 197.47015308582246, 211.6091200962555, 225.94200419111763, 239.3644792910658, 249.17334856554402, 254.47339070393787, 258.600071920737, 262.27110995300313, 264.4189542781736, 260.5566983655248, 256.573073824126, 250.17900237443516, 248.1571640118478, 248.36654689095533, 248.6570969983526, 248.82930075482616, 248.93143126800803, 248.9957861110171, 249.14832676081443, 249.26554137447485, NaN, NaN, 25.29193043587565, 25.436276566570783, 25.839207969638764, 26.387500457127636, 27.414203509934488, 28.369615375381372, 28.91633965644689, 29.8303301887229, 30.7096251626227, 32.288517519926096, 34.38442784078538, 37.43721831908197, 40.11727910404117, 44.161747443311114, 45.07614749710063, 45.552837524193734, 48.19494093419436, 51.76229767026951, 54.07832059504658, 55.43744857313853, 56.7968500247552, 58.921379345384324, 67.22293745821005, 71.33844890500477, 71.33337911063202, 64.93703592253078, 65.51576360598906, 67.7130615779665, 73.43652099217144, 77.62388020258528, 78.12574210794811, 80.53932701550595, 88.30418745997734, 96.3854814167237, 98.72294164438246, 101.79429581008877, 105.3230218090069, 108.62408480791376, 112.08587903878866, 115.91280188599981, 119.80064710870562, 126.7197315406321, 132.75741026037656, 140.7432801431691, 149.64026187892264, 159.4049913219207, 165.79410954296776, 170.54424024340946, 177.24163859412366, 179.75105755810011, 189.36117378502107, 196.9602034532241, 209.38557671128208, 226.378126647599, 240.59925093082458, 247.04416365448316, 252.75732487317785, 256.7673224769038, 261.40842765813534, 263.07668813668374, 261.0630511462874, 257.33970975859097, 252.5604880367636, 248.9595647417571, 248.56989340229984, 248.81617224645868, 249.00033685422287, 249.32748157572175, 249.35225485503491, 249.44397426660242, 249.61957761227308, 249.43861886136702, NaN, NaN, 26.54787631132624, 26.10201733820591, 26.61363860360701, 27.050433351026058, 26.973010505325515, 27.04203207659611, 28.58407439482271, 30.794764965581344, 32.92687010283123, 34.76216932681901, 36.964702470692615, 38.42828168121387, 40.85004810721311, 43.644565045073186, 44.234437836639025, 41.43305426641074, 43.26805931743352, 51.651107327222, 58.417065401953586, 59.739815726365975, 51.01643704743383, 46.665631922055624, 51.07120227974211, 56.87593932910791, 57.23830290096253, 61.13088176461704, 64.13360116399153, 68.89681390085107, 72.04618372304498, 72.11458735517166, 73.13000737666007, 75.39375875767051, 83.62220941774837, 91.03368527946618, 99.40085690791268, 105.35502859237249, 109.92557354918942, 115.37411724351887, 118.66869144158265, 121.46994935433206, 121.56075462659702, 125.98260596349165, 133.2639855929301, 144.73804492443463, 150.30355517763692, 158.0783346880274, 163.3737869349048, 173.9462911537061, 176.08164834819132, 186.81504982112992, 210.5854300754249, 215.97053631723446, 226.1780202753915, 233.21812451888755, 241.7979605565123, 250.24086008654328, 254.63762627147202, 260.13287932555625, 264.98273901647553, 265.9690585808068, 261.72414744018084, 257.5193584541691, 254.391028939696, 249.9061665589988, 249.2818561431462, 249.52185288097678, 249.8447385031828, 250.01469689375577, 250.10550668092816, 250.2130420384264, 250.33311938357713, NaN, NaN, 25.260580930295674, 24.81535723107449, 25.179344431967653, 26.2807043335477, 27.529522801910467, 29.809865672636352, 31.94122535328289, 33.62893003189261, 35.09836846113353, 35.97654069929478, 37.29934794425723, 36.41281568081115, 35.2290785776778, 37.8728863805472, 39.337559035856614, 39.99527774552196, 46.536840488856384, 55.139040533589366, 59.035826088668834, 51.83334402566457, 47.30185712595777, 45.38199762997657, 46.55068882998571, 48.45269929583195, 51.6763112061412, 56.078919165596254, 60.7868628542336, 62.69306613176841, 63.129205813425365, 63.71415446244231, 64.43645219204265, 64.4363013793461, 64.71736785385244, 70.8863558394049, 81.7649872892941, 97.48369653201986, 105.70759512705293, 108.3705189318722, 112.1981376374239, 120.12048687378616, 124.55619013653103, 128.76831044854438, 131.89812557889408, 140.0047434335552, 145.0018262639107, 145.8122464660295, 146.7631138725584, 154.30446684100562, 158.3853483806716, 166.37878376025753, 182.5128155206755, 203.12773442513102, 216.83198439199907, 225.76596908576826, 233.50446293558358, 240.599512966501, 246.660337059228, 254.2161160141926, 258.2984133326898, 262.1255068081129, 263.6283293988534, 265.77531654948103, 264.72558349906495, 258.28280926764387, 253.6826698611638, 249.2135900050899, 249.09287607674116, 249.34089265939082, 249.520273650807, 249.68927285610886, 249.86568516155276, 249.88443455189753, 249.92770902683836, NaN, NaN, 26.184071781814016, 25.810961311904787, 26.763665787521436, 28.45441536012877, 31.472335401932177, 32.12948481498033, 31.31557122741948, 31.458110710185554, 31.602387849563762, 32.04086772877239, 33.95245698942905, 37.77910944659805, 39.175708995173444, 43.36824214651903, 52.19620518380823, 56.24091636389677, 53.88783296645862, 48.58688464674295, 49.82860166696221, 55.192437221149724, 57.986880091646, 59.15468130358606, 59.00085597490061, 58.11945078968264, 60.17953290274318, 62.092785743613426, 61.79305542459421, 61.19635857926032, 62.069305711275256, 67.79834359132231, 69.99318519816931, 70.86696454175166, 81.7426018539226, 95.99753463636011, 98.33519059036395, 106.70853200540373, 108.03197621620306, 104.51020527642734, 100.09479472223677, 95.38932655041711, 93.436553307406, 93.21568378975992, 106.00866627727349, 121.89224670103843, 121.00153006498073, 121.21796095832795, 122.55635594334854, 123.67419285487017, 129.43130586456994, 138.5259418829157, 149.81842848362678, 167.16315230943601, 189.95265308158451, 216.06122852746282, 226.2725941656888, 233.34675839123992, 243.70789666166132, 250.06918074465457, 255.0192728662893, 260.1453931398989, 264.47865430045596, 266.39332709070743, 262.8722330362167, 254.5932315767152, 248.81158531251006, 248.348445407045, 248.67638044621484, 248.91995320178188, 249.09249936523136, 249.18796099383138, 249.28028662799835, 249.3748714717579, 249.42195402585298, NaN, NaN, 26.375201842524017, 26.963553715954408, 26.88669313965762, 28.430432640362977, 30.12243298330537, 30.707892639130584, 32.54668843894411, 36.37077557111482, 38.205020315283065, 41.29667959182936, 43.64937169797108, 47.03202036320535, 52.10265844522008, 55.55868240784596, 50.10949812472293, 48.03444922088364, 48.02367145770331, 49.044738658750425, 52.49934402383948, 56.471785700838225, 57.06197881500344, 58.382766326703404, 62.796321609909846, 70.18044103754343, 72.38372355688765, 65.2049157225826, 63.322445775538036, 65.74325857506305, 78.30611238966402, 91.09547835924171, 99.70188644697109, 95.86473269350714, 93.66631871231316, 90.78864556199558, 92.98471732989431, 98.60217813064777, 103.56729087754377, 105.88613128139389, 110.29357593656506, 112.7055767922831, 115.05672239877003, 117.39045415670054, 121.26881733568028, 124.87199825441367, 130.5675171137305, 141.94503566632665, 159.81769104848664, 179.8874327877044, 210.1058513081076, 223.67639017702683, 229.4930466480635, 232.90756545001702, 239.35913265755897, 245.45202391889492, 248.6568150105624, 254.91643880157824, 259.5314266056044, 264.5234397118514, 265.5758554268032, 259.10955615704484, 250.65616118179167, 248.26113138562155, 248.54331903981637, 248.78583125722295, 248.995431644047, 249.1379655294313, 249.2329787319012, 249.3010602209048, NaN, NaN, 28.524624760945606, 27.48660266823192, 27.702253080621276, 27.40175716386555, 28.871914136781605, 30.34003395138896, 32.76575449795707, 38.44065478363825, 42.045321773091814, 43.73255702081046, 46.080173970922985, 52.18738499325232, 54.16161583010626, 50.483428341476376, 47.82162576900876, 46.930093408636694, 47.28524363834449, 49.85336972537146, 53.969732645946884, 60.515631860199015, 60.77212543970899, 57.12196699641258, 66.60384060885269, 70.4694832336477, 64.9473074337667, 64.827706790094, 68.0140847182008, 72.41430374515141, 80.01826430865124, 89.3822451800162, 95.99269441571745, 96.99230947128926, 89.82359587256022, 89.71914208591919, 91.37580779244716, 89.92564784659959, 91.45339580479683, 100.05646686964103, 103.36503427176937, 106.11514447631004, 110.51439823233285, 112.93715013988793, 115.36741992759805, 119.36406828483975, 121.35847543974371, 129.35949295153534, 152.91247713864277, 170.2804004931087, 181.15802087820393, 194.06133331110146, 213.93572496365383, 225.9111767353512, 232.24559225156688, 239.27614354319613, 243.90720752900822, 251.2322750162173, 255.58490870225913, 259.0880441781199, 262.4028311656509, 264.77728029721624, 260.10604490679077, 250.31526602777848, 248.74121306429646, 248.90816900872565, 249.30235627939223, 249.36984127756907, 249.42874650863115, 249.49826889353932, NaN, NaN, 25.336733036364762, 26.88304468835589, 30.202427173981945, 27.917256211418334, 27.17239715180237, 27.45955114087259, 28.632590393657082, 32.31347604814368, 36.36082242925942, 40.18761279127388, 42.391070880237606, 45.84684493459398, 50.40040436835477, 55.83583052347555, 55.61206972656554, 48.40124988715214, 46.844759863161, 48.38040544366545, 50.50850253089235, 53.515249162792635, 55.16627642205707, 57.14644353299297, 57.2147713769451, 54.78287880004645, 59.77634957897204, 68.30395868726433, 66.53281367610255, 66.2273115881106, 71.43568302532744, 79.36780334015259, 87.81932267092077, 94.21608957951703, 93.4866863893261, 87.24027942758134, 87.02133291677465, 89.3734049893825, 90.39364987336643, 95.01517679273145, 102.50439983624412, 105.2336655313307, 109.32155793052799, 112.64192924163132, 116.17291627260033, 119.92233350580872, 120.35981978536094, 114.39720985850448, 125.25403316777482, 150.31984351777285, 172.36839551723867, 196.40529580709, 215.8113187841019, 227.17147424927686, 237.86004536841432, 242.50719180524396, 250.79356957297384, 256.9581740950406, 261.8373435727712, 264.50707949899373, 264.3173751165219, 263.6642380667257, 254.74471816243727, 250.0458915660735, 250.20686258724405, 250.52376584661528, 250.7612750612045, 250.8623558905093, 250.959230459194, 251.08014601835407, NaN, NaN, 26.14502415683362, 26.657711574765862, 29.752702302648885, 29.60548843910195, 27.390873628957607, 27.16245473505795, 27.893212693433753, 29.656244730509023, 32.81971393577872, 35.90781321230436, 39.66033240022343, 42.60253635060912, 47.67881466895665, 53.12111226420879, 52.3211233494489, 48.48408159741287, 47.51479188928648, 49.124867648823674, 50.587091898627605, 49.845865024289886, 49.32775553198909, 54.479188248721556, 57.0498268663009, 58.435820947835396, 66.73976993424256, 66.37357977997952, 67.16934090719279, 71.05922749924743, 73.2584856977764, 74.06032517419645, 79.93307543550104, 88.38844144369854, 86.552341587527, 80.15036456904924, 83.97883634694253, 87.94393680775791, 90.06087118947528, 93.07172545737284, 99.25272416076699, 101.82836158462896, 110.14040850313968, 111.02786115071471, 111.90037474630087, 115.85731352386847, 117.60408747820969, 118.47320907923566, 116.92810888818957, 111.64270002867462, 126.88011660087814, 151.30459835240592, 171.78881934859172, 198.52484004472768, 220.93948426161728, 234.80606526953878, 242.56837257125028, 248.5779982329011, 254.03742065371654, 258.461095594825, 262.70866453278404, 264.76280519270153, 265.17818750360607, 264.84278210750006, 260.81717471550775, 254.62160798932123, 250.12585944229247, 249.78485248481402, 249.81618818169298, 250.0535367588493, 250.16713020255213, NaN, NaN, 26.142538464020042, 25.62218999699626, 26.505915524501763, 29.597243164215673, 29.521501790607118, 27.454544929926367, 27.74382220757325, 29.581351314553633, 31.85773833586154, 36.27289502673607, 40.02472830449859, 42.375602391323945, 45.31647872976131, 53.41340699721835, 49.74111560160931, 47.67262393901346, 48.77077505230584, 49.871082316487914, 47.66378739470989, 49.134781033533365, 52.92409066661417, 56.818593501845875, 56.22297358642148, 63.28006885572088, 69.52374135242556, 69.7383597199135, 71.64219864705395, 71.27253695510376, 75.09253092448044, 76.20010031529974, 78.83616471988418, 79.57120516387481, 85.01528197435414, 87.43859442209276, 88.1517608772346, 89.09308081026293, 94.31197628572151, 99.7456014128999, 101.66319469555765, 106.95805673412802, 109.9008539873766, 110.12107491355503, 113.86275413830084, 116.93821434890349, 117.80550518272719, 114.49971237688641, 111.41791422137089, 130.44728936724155, 150.88891631309997, 168.25854773473503, 194.97189234544615, 214.79629314531965, 226.53983179988725, 230.52956258081926, 235.1408189915653, 244.4362810425255, 251.5138608000158, 254.68642655939357, 257.19554611494596, 260.99745546526395, 264.29371876754635, 264.50968006584816, 264.1224443073898, 263.7315433605716, 263.13715025826957, 258.771499391488, 252.5178949068316, 251.73956389881863, 251.56954251949125, 251.8893595395542, 251.93386672544023, NaN, NaN, 27.656462841558803, 28.31567584523367, 28.97477983089107, 29.707865840869864, 29.559160000574725, 31.471070471035286, 30.29001427813427, 30.062101695789405, 30.42093782404515, 32.69829732930233, 36.07857629919399, 38.13135708219461, 42.17981214374995, 44.7524966366233, 53.21278700931112, 52.85670018554499, 49.39082881064332, 50.341998820396235, 49.38256849208505, 48.11912600092063, 47.70485832980972, 51.523508771966156, 54.24244052871618, 57.69430404771514, 60.417044448510815, 66.14713308771444, 69.52346015296945, 71.35073978076942, 71.19249754653104, 70.08400847670427, 78.45479544102274, 82.78870305392627, 79.62665444633329, 83.3770161691193, 86.682064344557, 88.95273572835433, 92.47739801190887, 97.92314240621569, 105.78950752834632, 111.45414754459219, 112.71234829482303, 113.8083178645885, 115.34229147817709, 116.21425597953956, 113.3464697691129, 114.89494585388088, 124.61147774351998, 144.10267961779533, 158.8054812914272, 174.16243197007338, 201.04567975284263, 216.72384047283376, 219.62584315464477, 227.16893502817044, 242.908603214535, 249.97496002983095, 253.24124418696772, 257.5760981165106, 261.1978847645595, 263.2057363158796, 263.4658283107993, 263.3880770843726, 262.7969876396087, 257.91482918027145, 252.74494720514355, 251.82016236645126, 251.98231239636021, 252.32581890436117, NaN, NaN, 24.22607693110948, 25.18196075200939, 26.726476097875043, 26.35485306840534, 27.08922911644757, 28.929097575432255, 30.691727788409946, 30.026937582921477, 31.793006193928747, 34.8069366757992, 40.919484858039816, 43.34162969722423, 43.92038646323408, 45.16705899597697, 52.07981210558212, 59.28942491126813, 56.785871026120496, 51.40516140650765, 49.780977379893635, 49.47912726797981, 49.91428635872989, 52.33500470723772, 54.544000085634785, 56.85852888570666, 58.068383901067804, 59.612173852234285, 64.13275628781811, 70.7491361877595, 73.50364829790888, 71.72835867496876, 77.8925654645289, 89.12694670169252, 98.83563816556507, 87.48775641942566, 87.82229666299114, 88.13445402176636, 88.11715016979714, 89.6485078217044, 94.72771285855409, 102.68077953935374, 108.90382489935264, 113.66717545521065, 119.16634901765016, 118.9865982065788, 119.71666767587045, 120.63613141613402, 125.07108589431263, 134.1010467423847, 145.58093023378814, 161.53990560112973, 183.13687248940843, 205.41060571979003, 213.9735385072775, 215.4098669133659, 222.35102348732414, 235.40667067417624, 246.075623967136, 252.06452179151722, 257.6644030907056, 262.1460218544027, 263.99010509364643, 264.1682216738475, 264.0680863902612, 263.449823808586, 259.8717177565699, 253.3373643995916, 252.3460135905204, 252.66481733506677, 252.76528928056277, 253.18096355434417, NaN, NaN, 26.853028010899482, 27.291414603041368, 27.50978652321319, 29.71570440130117, 31.698235378127084, 32.577453527919715, 33.68082892595767, 35.22350436787768, 36.212613268842894, 38.08197656670742, 37.30408360112178, 37.95604884285448, 39.60721623670514, 40.264174065575624, 45.77534365433292, 57.25012682117401, 56.921762229040695, 52.83418534835231, 52.71217986093169, 53.140170990944604, 54.41220605747602, 56.49276287239014, 58.69780797961482, 60.897371283306335, 60.01163733629599, 62.32164248706019, 66.5080153471665, 77.64205104829045, 83.80644239037203, 93.6147531296434, 104.09680614062754, 99.14401453911385, 91.42833814682868, 89.87874155455575, 90.96141143308267, 94.15573561664038, 100.00369706373107, 108.06602180342581, 112.57476418518276, 114.9077981824693, 115.81341285585872, 120.60742590469337, 130.0096132082738, 141.08695909628977, 154.9758508976317, 169.2254112655649, 189.96423864768326, 205.79535472958864, 216.8617270913649, 225.7385757631245, 240.07582411195656, 248.11111797748617, 253.6691120390557, 257.7358354401678, 261.76377602027736, 262.9749545284158, 264.54363964321226, 264.46708081574485, 263.7219736663458, 262.9666561405128, 256.9916050968082, 253.36956899458457, 253.25480286956062, 253.35734687932916, 253.64214921830362, 253.66117111389616, 253.84242581929172, NaN, NaN, 23.96697483131655, 23.89003910957913, 24.477354445231256, 25.506191230228005, 26.901184895614865, 29.54876393697912, 31.384653743794107, 33.14558180129519, 34.68636869339689, 35.85889095256172, 36.66442014681849, 38.28040223046357, 41.21658371368227, 43.493428491811706, 45.991909824230426, 46.35541805476835, 43.631324268004484, 47.59572131620167, 55.607998971749176, 56.56654512641735, 50.42154817101768, 51.44467333287792, 58.05629929999922, 61.43483068953114, 62.974228234954936, 67.74977004169291, 65.90790158474151, 65.456956245275, 70.08316231408861, 77.13704248680268, 84.4047736668444, 89.75835036951288, 96.58526022683084, 102.38838933682752, 104.3009471879992, 102.26705422607986, 95.89027920968798, 95.59037538828518, 96.7003517105819, 97.42586875063795, 101.64162054528417, 109.8759487638304, 113.54403426794363, 117.38255388415831, 124.75385621421484, 138.01459628607387, 148.79660788660058, 159.7705768070378, 169.58448995411572, 180.24099126549658, 185.52871073344355, 199.18916884894327, 216.59993788489163, 233.77286885113293, 243.39179279006584, 247.05882278286467, 252.95068885117564, 256.21020245814964, 260.79848423572025, 262.84976695630974, 263.7068990183462, 263.36200705428564, 264.47666911381066, 260.38594550923847, 254.33263977190973, 252.53196777579336, 252.563463749937, 252.7395454627312, 252.90829948243402, 253.00336103489053, NaN, NaN, 21.195670453405842, 22.188916135029366, 23.84468442553567, 24.982391042121947, 26.08621539824771, 28.18082807625182, 29.243930291938494, 30.303790313269573, 31.143566906352177, 31.468935625804686, 32.89726479083633, 35.13542182624413, 37.115381996247535, 39.31703077430115, 41.81761420101114, 44.20281224264166, 46.99730677916215, 49.96946302093443, 51.9870405951668, 55.2596482209395, 55.36208942901638, 55.46401849150705, 60.41453325871219, 65.37141434995536, 61.95170812300536, 63.70954631779747, 63.70202712346572, 70.08734640163122, 72.84437483412111, 74.60728879080663, 81.65851432914495, 91.24039985812924, 97.62232222031535, 103.67878044041737, 109.19663028359317, 108.65982730615914, 113.1896717710949, 124.2245417525078, 126.56766350088466, 118.30581753648873, 123.31909364748486, 129.3658165421984, 134.5273628158968, 138.09117488120597, 145.7971191633128, 154.41286434922225, 168.69095213859794, 178.77205266829776, 196.62490287706288, 212.23765730759553, 227.9582624610713, 235.25937655620092, 239.5139578370475, 245.29373348512348, 249.44183520468562, 253.75132641167102, 256.7873980184183, 260.6507780103785, 261.7313348623411, 263.21850296252575, 264.0170144793085, 264.8415017786221, 264.6063162137331, 261.4610937242732, 253.97059248816254, 252.74138143019889, 253.06719810840985, 253.08621366281625, 253.28233864447057, NaN, NaN, 24.372857063040257, 24.370270771466448, 25.510779063415836, 26.280719230619937, 26.717963932115318, 27.967499951129707, 29.40057940757987, 31.681505668347555, 32.34289900608085, 34.291992817844246, 36.42653351390093, 38.29715581578848, 39.72668157276916, 42.04315249436061, 44.72656812848452, 47.25858769793706, 49.82988165785655, 52.36181768922954, 55.33108981986331, 59.109793823587864, 62.37292959399333, 63.47006330704947, 64.71290343406612, 66.98057955294188, 71.24018558438254, 74.32412844237798, 75.34670531876223, 72.4035660344671, 74.14975721474285, 75.68078948753491, 75.006689710218, 75.43666739083406, 78.88213121022946, 86.43556894654806, 93.33864312987546, 97.74245057890901, 95.6870925616293, 96.42152337905047, 103.98245416334774, 106.4886356356988, 106.87554642117236, 111.72726519645916, 119.54310237853859, 125.60646892608379, 127.55592930776105, 128.47265078117093, 135.588865493972, 143.86130592053925, 161.34492375945868, 174.26994523538778, 187.32686087168622, 198.08252238221925, 211.58201605490737, 225.40249765356623, 234.30238465880825, 241.34738963537995, 246.3832333376551, 252.03894626742203, 256.95891715961295, 261.49541718795825, 263.3507381790049, 263.1634448406584, 263.4037000126485, 261.99988175571747, 254.82818832662417, 252.1294389335514, 251.588101873147, 251.8327900437963, 252.07658316244923, 254.19743254436182, 255.25868899054007, 255.13073800330736, NaN, NaN, 253.7922838423942, 253.81747895562583, 253.84600804228634, 253.94078409694833, 253.94548179696878, 253.91521861049827, 253.923978697337, 254.01662736956325, 254.0840723573345, 252.91748258968482, 252.97496754136924, 253.40224075349477, 252.51708363892004, 252.579545295633, 252.45651352564414, 251.3347422480356, 251.565538102904, 216.6177812243208, 86.31386081935419, 61.58153836564415, 61.86084428637735, 65.74674464664233, 67.87087175894517, 69.33296964204763, 70.65639167776595, 73.88403641581742, 75.4848901247146, 77.2442953546329, 79.58584219048734, 82.88937080849597, 89.3353141230066, 94.76540462325362, 97.62564480952453, 99.39641974987522, 101.1576299358205, 104.0252502140031, 105.72447978051454, 105.89093163436402, 108.61953236752805, 113.10802345082419, 117.91919047976906, 128.03464775492657, 134.31978813936738, 141.3408495412661, 152.65231724041297, 169.4671256937398, 188.61437302860085, 200.7147427449083, 214.34154060052515, 224.6470242484939, 233.6891998403054, 242.7556271215318, 248.11908906401763, 251.48337881583595, 255.37795250414203, 259.4721820042675, 263.4726950631407, 264.4915238799946, 264.2257173362035, 256.24306423658044, 251.7958268711613, 251.36255878922748, 251.08657439801271, 250.76358529824083, 249.5340417664957, 249.1711959739924, 249.09940690996632, NaN, NaN, 24.922106606522696, 24.660119939866824, 24.72828509375323, 25.274414359102604, 25.709881377251087, 25.854047729663957, 26.88144011994814, 28.718020740999798, 29.116807030379434, 29.075104263751516, 30.097848198111826, 33.477765546969856, 37.00638967468955, 37.95784538359949, 38.42730649841856, 40.443371124691296, 44.33408760048329, 47.85819547096147, 50.67976876654289, 52.51220598737166, 52.063516288223596, 54.47962596895989, 60.4267706143667, 64.72501119910571, 67.3665723992014, 68.35238318106546, 69.22632788113887, 71.53694836756408, 73.52215750713286, 78.03288100225218, 79.35920262168139, 79.7903175553585, 80.33239277368149, 82.5319838393803, 85.836345010112, 88.80574928031058, 85.17578320681008, 83.19424927206282, 84.28600335222474, 96.28941424574691, 104.90548006776137, 110.37072277928185, 113.46606237276644, 124.21958190865891, 136.0221392910882, 143.26483442810496, 154.6496932559512, 165.78197555295068, 176.37253413166795, 185.49249073621934, 198.50651516669356, 214.6877017118266, 225.9509819433698, 236.01823343835272, 242.82772422762136, 248.9951445374831, 253.89641668828907, 256.5030070735777, 259.9323107720957, 263.3443531607177, 265.4930002322465, 265.50547890813004, 261.89182564580057, 252.96619544903388, 250.65531502328952, 250.84808391667227, 250.83042045731574, 250.0557267444252, 248.6783212604824, 248.64916094769035, NaN, NaN, 22.149384972008352, 22.296086300248813, 22.846643859023562, 23.872899380411447, 24.863950253501127, 27.625076447755667, 29.867948901625887, 31.18662168368748, 31.992568746594102, 33.49924938798738, 35.259901011594245, 37.16390049167275, 38.95718635015479, 39.20875388815881, 39.753858173035454, 44.01543368689123, 47.65990012473, 49.34762141308156, 51.287128178242114, 54.95450512247823, 58.03298564832189, 59.89799248829779, 62.20543246936147, 64.18871707667057, 65.29027932768835, 67.82965098521764, 71.58276603187147, 78.40922064454232, 82.70191918530826, 83.91623493262043, 85.90465439682771, 82.26011334819978, 84.00499129884301, 91.26540377987641, 94.79755085039213, 90.06234776608304, 90.7228131852584, 91.70549360873414, 98.42317796176263, 109.55054645173622, 113.86494117093417, 116.38047222177087, 116.84416813086527, 130.71675706778024, 143.26519364270086, 153.48914423643916, 168.93371055764408, 178.77672318881432, 188.31542897554567, 199.04359451357175, 211.47533977590396, 226.87858634168447, 238.25037363774624, 248.21892095925045, 251.492424069995, 255.79844566373376, 259.47439364590326, 262.29103776355873, 264.09397730784116, 266.0862273364447, 266.9851292441303, 260.58747860105984, 252.3501414578397, 251.57210156085318, 250.55045400478016, 249.86689594827055, 248.02442073311136, 246.48339395522353, 246.18053636838138, 246.5381472628425, NaN, NaN, 23.48784600631909, 23.5584175491109, 23.959601293150353, 25.022559918334288, 26.934282325414085, 29.285466896801577, 30.936933725148307, 32.44007136892288, 34.200617130727224, 35.81269254680137, 36.91013511797521, 36.978886140299366, 38.81114735609731, 41.014198547761445, 43.25217331838855, 45.5650194411642, 49.047287199177596, 50.547547322219884, 51.785253430912995, 55.196759459846106, 56.368063534964556, 58.49492122188108, 66.6424974676999, 70.76444934554063, 70.39797620584591, 70.83314643584458, 73.24559879696801, 77.71944261023148, 81.60630381762904, 81.9763078816847, 79.32932778792511, 77.64072842267787, 83.72280360377773, 86.36645937461056, 89.16058698284071, 93.34307951417581, 101.20746339373521, 103.65484191767139, 107.10105563106, 109.59304000093971, 113.37888715933346, 121.78682163711245, 134.22036354759447, 143.72640264482803, 154.26856435741067, 170.45811384056785, 187.29373436487546, 196.1866645749562, 214.27008078489675, 230.40566702417865, 241.55290895427817, 248.77300716655904, 254.28460721255857, 258.9195090674149, 263.7913146534133, 266.32097842658, 268.03655406201847, 267.418608037344, 261.8176500180895, 253.36929627738024, 250.59065186659652, 248.7244101304013, 247.6238900302599, 246.90316787520226, 246.51680291439493, 246.27171529430217, 245.97987825415808, NaN, NaN, 21.558805085169517, 21.482929647148413, 21.737933939148114, 22.507961183555707, 23.351388696272632, 25.668998901033216, 28.648776973191154, 31.62438710036343, 33.90256787329612, 34.89255133256194, 35.40288588098103, 36.610354901610144, 38.07536572476554, 39.02581873392504, 39.39165786069952, 40.45337433848972, 43.062812158070734, 47.03617445975762, 50.818320583978256, 53.901696500515804, 58.013573151548826, 61.462644287542965, 60.206491072494636, 58.28997140741683, 62.32896967144364, 69.599613216701, 71.21774805493676, 72.31966469618224, 74.59254827307798, 76.19584503976508, 79.86135507233533, 85.31211771189999, 84.51936151302277, 81.57560436940285, 83.62402800318672, 85.67001849277949, 89.48126489954919, 88.58670432275588, 90.48295323849099, 98.49000243756578, 100.0071081358469, 105.52977078073691, 113.44020517692184, 117.86184348832136, 128.93202853023092, 138.73261678657593, 147.7719794944494, 154.9862613879334, 160.05278279525496, 168.61273745171187, 178.28970939151267, 192.99710725271012, 204.7149850624625, 224.8423675195162, 238.77300944300157, 245.50840437219702, 249.85554637457753, 254.49000845869566, 258.6723480008297, 262.1512689948434, 266.88506085235605, 267.77543434063836, 261.0617280290614, 253.74935329681102, 249.49062894198843, 248.96871635361305, 249.44206946090347, 249.34853363169134, 248.84052178609983, 247.60465903358946, 247.17184282107067, NaN, NaN, 21.303711350666205, 21.33775956932482, 21.887092633765374, 23.35694355873693, 24.824756615240325, 27.43243991944322, 30.37420620200196, 31.839554384243275, 33.30872285639525, 34.63214538622534, 35.548809700198746, 36.390663325533424, 37.081844115758415, 38.105087996601995, 40.162890874888454, 41.5557524057735, 42.06741072023655, 43.46111753802166, 45.294303964432, 47.97228042803912, 50.17668635584313, 53.18293591966205, 58.61043683730525, 63.00780359521036, 64.7652426682247, 68.0667089993597, 65.79403743359683, 69.08814469850753, 71.95217385030493, 73.3468914960999, 74.29984466599531, 77.38211087076412, 80.31008980589759, 85.07796061207537, 90.3635639776416, 91.98580559050536, 87.42739692863508, 87.19894797468709, 91.52811055029838, 95.56746839132263, 96.14972247960293, 104.51511929519108, 108.47973432556661, 111.12585729142769, 115.09528346789656, 118.07707764687504, 122.17878363627192, 124.22403667918528, 131.6543302922779, 144.84124635564942, 150.86315939868166, 163.8855688691145, 177.49551586080972, 189.1039348788173, 199.71632524657204, 205.2815277002312, 211.7936054408003, 219.82810280305907, 230.1034953511598, 238.80800030230247, 243.8177793121005, 248.88526495352545, 254.8785681538595, 260.6527807948851, 262.66400896538113, 262.5356959556318, 259.9411316688745, 251.81985915441928, 249.10166821696367, 249.34696404561026, 249.60279491475262, 249.64278545995109, 249.09367928911777, NaN, NaN, 22.924291215877044, 22.2954986257626, 22.623017891066453, 25.56416756665099, 29.499803815722803, 32.072677786245535, 32.98714042427955, 32.8339445731035, 33.49259818970274, 33.891024304951685, 35.98367129014639, 37.96277590894452, 39.428876347090636, 41.81398203531724, 43.13458598022031, 44.45411327039092, 46.47099406064557, 48.41399282369985, 52.59786903094238, 55.56915830144296, 59.381962854933, 65.32918405619307, 68.96118243800049, 70.38656515331851, 69.167598907388, 67.61926464338575, 73.33928680760398, 78.19409549875898, 81.9442048031078, 83.92580327289825, 84.35315632960388, 86.32754635006883, 92.50673018128607, 93.05537238449057, 94.48634781824907, 94.93283490351148, 99.55142033238361, 100.20291448481429, 96.24353915938228, 107.71068157347537, 117.31765517069717, 122.05234873296021, 121.93589761519324, 127.85825789175274, 141.75417135800035, 150.3958333633047, 164.44420916170958, 175.1412619040059, 183.9001240043914, 193.59607302887963, 202.55782698410997, 213.49684744397746, 222.22757681863865, 231.43810624186048, 240.71042231349483, 245.99125290527547, 248.9851683971997, 251.7952363503293, 258.24085648605796, 261.1303789882261, 262.82192198847315, 263.94003487192805, 262.4767115575069, 252.47229985449658, 249.58936549096703, 249.44369372734042, 249.41020622144887, 249.05827868092518, 248.11553719810274, 247.89491858395857, NaN, NaN, 25.652841532401624, 25.206326012576746, 26.455131705447098, 28.36563643502997, 29.98246568910988, 31.15508896483024, 32.03253223120575, 33.09293798691342, 34.15643495956283, 35.36405124884207, 35.94636317840649, 35.94104421435955, 37.51588376770436, 39.420770249279514, 41.327169937942706, 43.26994786958847, 43.592225064792345, 44.17443953574209, 46.78206542660271, 49.45625366349167, 51.40176799606656, 53.30657372876148, 57.85056131416775, 64.38320308549328, 69.44200659062275, 73.47564570759249, 71.63853276715965, 71.56429855499582, 75.31618059647151, 83.01924637988897, 87.6429946308429, 88.75644985046935, 90.67070122900316, 93.30305511595235, 95.28891969266365, 96.98112961951922, 99.19138603577906, 100.22917039334077, 105.00885826047742, 110.89772849685595, 110.21941677827024, 122.52655100526617, 142.97930457744368, 151.92232663947408, 162.29253548018534, 175.71045083797654, 191.52280495832497, 205.90669099007525, 216.57797432574304, 229.03136084538193, 239.44029780517556, 245.54633375945, 249.91466538453872, 254.9929271562293, 262.2867121601881, 265.57616353045364, 264.56496807696107, 263.3008172165738, 261.6562560699711, 260.10092550766234, 256.2453106408829, 254.03231485209483, 252.0599256726362, 249.3484359787459, 248.07596120426058, 248.18718068457403, 248.41912149891667, NaN, NaN, 24.39443915664378, 23.83793795939749, 24.75645701910413, 26.48292507683478, 28.2096449431594, 29.863224908564554, 32.21627997061758, 33.24491383418324, 33.828249775735344, 35.07498487835386, 35.328720362076055, 36.27844062308614, 38.47769068913537, 40.05193013607993, 42.031754141963695, 43.45480206300818, 43.37215004560782, 44.172380976896925, 45.45002544193958, 47.79487772015818, 50.87592767791967, 53.51638618130603, 56.07734524481222, 59.22895560623408, 64.94863929503592, 69.12876938315902, 72.1369039522421, 70.3002047444545, 66.10708402704192, 68.5292396335672, 71.17004575743836, 74.68217423966868, 81.20323015509595, 85.53251294985971, 87.14424558591163, 90.52877755055128, 93.39004892223606, 94.27558922971645, 96.61956983502064, 99.27451196225049, 102.1531360994222, 106.02841306359558, 108.98688500788533, 116.00311175558905, 137.16000781997298, 151.606919738498, 164.67141702847445, 186.82262576168378, 203.61589651286877, 213.0546257457534, 219.82550987947567, 228.08888115627119, 237.32410750859034, 243.79613579509896, 249.0950087539343, 253.32986808960212, 258.3844841424484, 262.6070564335954, 264.06769870237844, 263.6732272553881, 262.69192417664215, 260.840985037835, 257.3022323512535, 252.84926774487462, 250.91450794971507, 250.37970114274964, 250.24922832690802, 250.42868382812628, NaN, NaN, 25.870775190580165, 25.61027627552401, 26.084526543163136, 26.41065761282741, 26.184499193271705, 27.909794398975183, 28.898186818908695, 31.43542044255447, 32.39156476449624, 33.08542355557211, 34.589695581581374, 36.75629407499566, 38.958092779202865, 41.34240903338128, 43.21309280706205, 44.60776862585186, 46.03561123836557, 47.830303462714795, 50.57991235712032, 52.70351204812094, 53.50050339299118, 55.25231916612455, 59.06267361264662, 64.56068050241304, 69.10854667389148, 71.83299226457656, 69.91194816249664, 69.75375129886274, 69.89347254819715, 70.4792393776912, 75.0193947726804, 77.58353979580754, 83.74665660550767, 87.0492963138433, 90.13720287445227, 95.64901345083065, 96.89750527046135, 99.85771125076072, 97.75056807698688, 98.33507227700994, 105.42804340773995, 107.21356224056031, 118.69443386899866, 135.7767605200206, 150.6964459431458, 157.0875406097836, 165.91229761442438, 183.48233728161884, 199.12013017034164, 210.08996794314152, 219.29315493965737, 228.44852786502568, 235.1868933990256, 239.03360589678607, 245.45714922704204, 250.4671419917587, 255.30376062275582, 258.03282461228974, 260.3885082288746, 263.6998922598336, 264.3651716012192, 265.1578302888916, 264.6641952673486, 261.7055063163389, 256.3466794653368, 253.21326076837627, 250.52082587832092, 249.91749939502452, 249.82973892722484, NaN, NaN, 24.06048202797541, 21.62606452724144, 20.59097679389164, 21.323826746638336, 22.71940207456684, 23.96646477352765, 25.656537241745156, 26.314935727339098, 27.563208235240516, 28.956875790774287, 30.8645434051679, 32.846866348545014, 33.652560196814434, 35.0474221733259, 37.39774621951811, 42.09848798311983, 43.786547597146104, 45.400923048383646, 47.52855404006613, 50.82844523728666, 51.92440464204934, 53.685052002946456, 55.953045933678574, 63.953735602762954, 68.50930038957291, 71.23346759230179, 72.39723357676633, 71.44000364556778, 70.55514654800504, 70.77128262258128, 75.61478530563907, 81.1929136359639, 84.4200411576779, 89.0372812265571, 91.07832379764324, 93.50062669238886, 95.25212712492696, 98.64097326960899, 100.56039855197058, 100.11897163653256, 101.29847004085859, 94.9959139669918, 98.5030688809473, 106.73063499661889, 110.39690111276609, 124.41586936409105, 140.19782997557505, 155.44683220996805, 164.95729010535544, 175.25894688975924, 190.88058464006346, 204.16596099620222, 210.96298875520975, 220.56796005275825, 229.88538292764017, 236.18655886795418, 239.24559382536393, 246.09827742870002, 251.10763141649045, 254.25880313136406, 255.8940261993349, 260.0221358817254, 262.81802655436144, 264.48117472407864, 265.0549914257371, 264.5506749763318, 263.49583654650553, 255.88761243159743, 250.58070711663473, 249.82190071102448, 250.1366970659754, 250.25103172917932, NaN, NaN, 19.157434829515488, 19.007121432430697, 20.698682968966345, 21.72584862234667, 21.571180700901262, 22.15426928604878, 23.916889297863843, 25.975514198683758, 27.592059309337245, 28.542780822956516, 30.374897749768156, 32.064042743722176, 33.23717997598079, 37.57164721990669, 42.56709016161002, 45.067246065551174, 47.12144606815711, 47.928536025203414, 50.78556126551974, 54.89520996945702, 56.98292968938007, 61.38257430165334, 65.19770035086616, 67.83110564033787, 71.20659911218104, 72.80899344064717, 73.75772520605578, 76.03149997870757, 73.53634581849289, 78.81665276762175, 86.74222108683095, 90.85332661983028, 93.26624711254607, 95.69331937604113, 101.29546344029826, 104.6739537688777, 103.21290070147822, 101.31454584921964, 99.70551530696302, 108.82303824248109, 114.64006514741794, 117.29434537814149, 126.74825916453965, 136.92695285616588, 153.024432150888, 164.27757287768554, 171.89011545049695, 184.55721982511972, 197.7627792351771, 209.44714879883742, 223.9336666342261, 232.0223913200024, 240.17178778648056, 245.4002055995207, 247.37086480876206, 248.45778234048356, 253.6207805860712, 256.8013399397391, 259.7238663485176, 262.1241001975999, 262.6571937095781, 262.91446116634626, 262.54382050287273, 258.8954159027256, 252.89231824797633, 250.34764423646857, 249.74444061228482, 249.91827787317658, 250.02169653834437, 250.14190206234107, NaN, NaN, 19.560556519126795, 19.18971312907147, 19.73848255684189, 21.206902482706163, 21.573128332582503, 22.267302234453005, 23.32978797076494, 24.57596392634873, 25.491092581126406, 26.000311335011858, 27.134783557717494, 29.411855478183348, 30.91793442466482, 33.156690990500785, 36.425743695456525, 38.36798609296721, 40.67912094958336, 43.0667165761046, 45.81763563493848, 48.018469356808666, 49.89161154064356, 51.43384283317056, 57.04613676403616, 63.543750274626795, 67.3921357480692, 71.13139665577246, 72.56427542033748, 75.53206360937959, 78.38730653332964, 80.46974009053919, 83.88281239328093, 85.96907739163952, 94.88836211322862, 102.59422255019098, 107.86852350230504, 112.70451897770343, 124.70287960172449, 128.66046734340043, 130.1898596810392, 132.82491892339286, 119.00546473332706, 109.92204522165245, 121.68834586126651, 127.76058162857144, 137.79326821189332, 143.256430219739, 154.787399203126, 163.9880877673297, 174.18242483028905, 190.67090820944696, 204.59292388951954, 212.53338886633193, 218.96729195929655, 234.04857734336437, 244.6049571142893, 247.19847968318444, 254.38270004668988, 257.8788289457661, 261.18422327216655, 262.83969054222354, 264.01199737796964, 263.27741378169753, 256.1053884596102, 251.53924893711692, 250.49194632655153, 250.53193319301946, 250.35424730794517, 250.2572081628754, 250.67477787968866, 250.80111928496865, NaN, NaN, 22.624691872554713, 22.3643122996152, 22.546783285814122, 23.021764246479954, 22.870216530897423, 25.847295743174275, 27.428502238878156, 28.78388949293049, 29.992755070201703, 30.867980450815345, 32.51588159948183, 34.535156467643844, 36.11115348068115, 37.94294319921429, 39.587134985067664, 41.01042434967362, 42.764180622829784, 44.337897737914446, 45.363485286700886, 46.569707047354775, 48.692873608095766, 51.259530439566355, 55.47300319895375, 60.05508811559973, 65.37362267413434, 68.30850930345642, 70.69200691369939, 72.52413829933879, 77.28815890671991, 81.13548382040183, 84.07395601517413, 84.80306148176354, 87.73101771729277, 92.85839329067332, 105.33202391852318, 125.70200962114743, 127.72549428600657, 132.871578963824, 138.21045277257303, 138.79253373519398, 143.2050043748133, 146.91750451963017, 148.4465097909897, 160.49339956460187, 167.2907687433464, 182.63691510690853, 200.369188670614, 208.43725975328272, 212.62259150439976, 218.1021840964203, 224.7338832418125, 236.36462176321874, 244.23099815342366, 248.83282897494786, 252.92458437775358, 257.78955230350033, 260.20385631574055, 262.62120770817046, 265.90735969682925, 262.8183666647025, 256.6403519752979, 252.62887803005802, 252.18597563612119, 252.51791436046338, 252.28151763719382, 250.99268165479413, 250.2744650727306, 250.17185083862626, NaN, NaN, 19.34242161067406, 18.67548980228674, 19.335571519475774, 20.3611167248754, 21.240902583796476, 23.408783609944447, 24.987027569469245, 25.458766584308005, 26.85224880650009, 28.246676947666288, 29.602585692433845, 31.36229272094917, 33.673747422006464, 34.552021814180534, 35.43161283352408, 37.67088079583915, 40.018429194335475, 41.4467509257081, 42.72623752052706, 43.421544181393514, 46.20974205184107, 48.707171641868435, 50.02697362385507, 52.81138341452128, 56.32682494482276, 61.76004626066388, 64.98926979096612, 68.94723212073171, 70.12452038657456, 74.81472861922605, 77.8912275835205, 77.88572853854498, 86.53729356797373, 96.06904169651676, 97.8181045429873, 99.57583724187413, 102.94630262743226, 121.29671666195392, 132.01213787365958, 135.7003978469124, 137.9318654539921, 140.13959696645355, 145.48166334040062, 152.04664251827822, 159.14735247802412, 165.24724267202703, 164.0492406093271, 170.05356200247428, 187.41628905060446, 200.60699483943884, 212.971284224856, 222.0522491050599, 232.1302117590013, 240.4893077151506, 248.87580471046513, 251.96813501222064, 256.4799525294947, 259.83175778202326, 261.6327751877788, 263.3379613603419, 263.67328310166334, 263.36858221061283, 264.5924116681447, 256.467503922968, 251.96794457328528, 251.83970334016894, 251.68090488550547, 249.9151366429619, 249.96788110296052, 249.69649180977936, 249.74317313379234, NaN, NaN, 20.5966853093035, 20.48501989861727, 21.329174200534307, 23.13007593913606, 25.004953552047326, 25.259131044196955, 25.549525360549058, 25.80321468197792, 27.123180544903597, 30.208257695577952, 33.15013948229478, 34.14055047696935, 35.24291237434092, 36.673515745918245, 38.36292074659276, 41.40788024235465, 43.0943341676868, 44.22938532827009, 46.54663136822482, 49.4123135668678, 51.019865101762626, 52.48122780828852, 54.67810029093905, 56.13812439091596, 58.18517831139519, 61.40595911954247, 63.903027239715655, 67.8635112486677, 74.31163799254954, 71.94797835608534, 73.11181398737887, 80.88146392174946, 89.38560718053544, 92.02867204556684, 95.25832507032267, 101.99931819799482, 109.4822251942942, 125.76573529544869, 130.74541372979397, 132.93390548005772, 134.32186823201238, 139.9587946807935, 141.07676516482778, 145.75110208692314, 149.43750969011492, 156.24072402061893, 163.5929488902221, 167.56543202100994, 171.6999534183341, 183.95445309709692, 197.8118417928389, 210.82606271683713, 219.54104753845724, 227.24510900122021, 234.03458161239178, 242.76117314965325, 249.5070344279796, 253.31756880794006, 256.17629595409835, 258.4797124114629, 261.0576180610697, 261.95188181072257, 261.0527820271208, 260.7706034017282, 254.05017576798352, 251.0242374611186, 250.01513794926436, 249.29606281687728, 249.03226714698005, 249.20129602361737, 249.46416732101284, NaN, NaN, 18.93671116874204, 18.45492710128725, 18.783076192793562, 19.58896744720124, 21.0229052741826, 23.191767167139798, 24.880761408715955, 27.9687323863883, 30.026603190152148, 31.49022481636884, 32.33043737147582, 32.655735936089044, 33.49389112356622, 34.44716539198104, 35.47342943678119, 38.554598796086786, 41.96742991708265, 44.61266094348403, 47.0323920356834, 49.416388403747774, 51.249525076236225, 55.64757631852227, 59.16352738930709, 63.67008233665071, 68.73618076116423, 74.01759226923548, 75.00590803080163, 76.20934267112465, 79.39488854283604, 83.24305578025368, 86.43241383556278, 98.87105356505434, 110.20811196156934, 115.3788447072751, 127.2625902838272, 132.20971451045648, 135.07996203554353, 137.1832168519757, 137.32202768901064, 138.94852277117693, 144.0190674641931, 147.10880900171156, 150.95331127720678, 155.53494595660868, 160.42372884459715, 165.5733069103404, 173.4045488490091, 186.95058351537813, 201.47643358566003, 212.93571527144064, 222.3418550253303, 231.26356662801064, 239.97828426642837, 243.69049372519007, 249.66008044131158, 255.6632181832309, 259.7043932303926, 260.8639922310214, 261.2365358670281, 260.83261319099296, 259.6570997877839, 255.33100652860898, 251.64106408369415, 250.67769785381768, 249.61869148081746, 248.81037799118354, 248.47568105928104, 248.65582286705043, NaN, NaN, 21.031730469013816, 20.882593576906977, 21.3217144145147, 22.935940854731157, 22.270765773323948, 21.531040520292112, 23.00123092421528, 24.101302693242847, 25.421572695401277, 26.6687078231062, 27.325855039040253, 28.49795608683416, 30.478674588881294, 33.04670429114651, 35.68559909920097, 38.47412204177813, 43.173687303903066, 45.962430668473516, 49.11590023988438, 51.393145115482575, 56.78584691211339, 61.95657727152187, 68.89167577244689, 75.59829310640833, 76.91075129030686, 76.90183566134195, 76.24040221431287, 75.90853283476369, 76.67307469782924, 76.66383936313764, 78.96946099368037, 84.36044648973032, 97.77442115340111, 97.99156983771242, 98.53017510297529, 97.20331802737392, 106.77361352440523, 118.9853859571407, 126.34408737873778, 129.41116121767544, 130.23549519204573, 129.83546316484416, 134.10541451245516, 140.30778480496758, 154.62991655175017, 161.04376930599764, 167.96044289581093, 176.0294538844841, 183.24107809847484, 192.44680931835936, 208.06643372947235, 218.23464387282837, 226.15942411536832, 235.24283618881938, 244.12865621028547, 247.96001142346213, 251.8943143831588, 257.41161928186597, 261.3487320716195, 261.919386010618, 261.75829054303074, 260.75030522480574, 257.79207304608616, 256.18798275769024, 252.8699026001538, 251.14836653765556, 250.62213114186264, 248.75111803084573, 248.10225594179494, 248.05248313955903, 248.08106808084395, NaN, NaN, 33.44920139074846, 34.034752240321815, 36.16472645049623, 37.554656394224146, 35.48735513758132, 34.52137579382864, 35.470238381452084, 35.31615934681374, 34.647967575032126, 35.080975054051194, 38.01414882748278, 39.625505567168474, 41.09222973420167, 43.88183318097942, 46.010264905040685, 51.87969608758476, 56.871589460670066, 60.902782286491004, 65.08482599277902, 70.73751789359305, 76.61045194464383, 79.84231049627103, 77.64283565542782, 79.3246017922321, 85.55667882405295, 92.82880935917488, 98.47748422277935, 103.08909762302592, 102.71942896978304, 99.55553371229072, 98.21850624939816, 99.7454600242069, 100.53979771478603, 107.9346321788518, 111.3846981636737, 117.97540013301733, 123.84565087389473, 124.52262629808003, 130.11794431187795, 135.04547710636913, 137.16004081408659, 143.14533947903033, 155.30725968864039, 161.51788172526966, 164.76273483290583, 169.67234194374214, 178.7502884750734, 190.76723011205544, 201.09645292557727, 208.39682568431846, 215.54871428191163, 223.75215576305536, 232.1197537201496, 241.13957877112495, 249.69441434772727, 255.33546998463433, 258.89102341934756, 261.4913683344701, 262.4908008733524, 263.75597913634044, 262.64625544192467, 257.3671708091698, 251.15838695046645, 250.38400101704664, 249.59610458741918, 248.03656336791497, 247.1470751356986, 246.81667488087976, 246.77332959840209, NaN, NaN, 37.389424355922515, 36.97971151425478, 37.30850365306777, 37.893922742026874, 39.06665721541723, 38.9848870721641, 41.366565677275126, 42.53423497608232, 44.10765006669024, 47.19380977466106, 47.224921400932175, 46.74050405771351, 48.16880843803298, 51.726678667031585, 55.134611250853524, 57.99235304972606, 61.8820401201124, 66.32570976708404, 69.03740901011092, 71.15756352161769, 75.19422809284154, 81.49864312467135, 82.15071545134269, 81.19165684529258, 85.59825862275662, 88.67251935248107, 89.25420325816808, 95.26394072037395, 98.11785733054602, 101.49199062533373, 105.82122404105765, 108.7493266169716, 111.45768058685007, 113.94053475094815, 117.52431357333737, 120.24716939979052, 123.31310675884768, 124.11941749093211, 127.80017273620513, 132.3503028185984, 134.15399649705628, 141.64647392744948, 149.9055848869901, 155.68209017801482, 161.1815152075931, 171.22312500252718, 178.72620037773174, 185.34107637696752, 194.84253756666894, 207.05640272043647, 216.99422588754123, 222.3743288813829, 227.38108935992474, 238.26900333499094, 248.9304807972944, 253.43140114361853, 256.59135636876255, 260.42686442665314, 263.2085207543166, 262.47376806312644, 259.3061734743552, 252.9180219903419, 250.65613217559647, 248.83341544746645, 247.4083046479814, 246.31756236424584, 245.99044012542737, 246.0927454384025, 246.26589890791135, 246.21929280320808, NaN, NaN, 35.18514337395562, 35.989918770251954, 36.0617189323603, 35.39217079977212, 35.67979017764722, 39.353805753508574, 40.96719697189251, 42.06220424093983, 46.24340344173907, 48.73651228671291, 48.803683462241345, 50.927369720856525, 52.756229722769014, 54.36391787013704, 59.35479170244137, 62.28496831333306, 66.4667541553505, 70.13318345873355, 72.26148499357103, 75.11469745329322, 77.6354602144198, 82.32904196984579, 82.46378169574453, 85.16806538024149, 89.48726353994068, 92.05770935264094, 91.3181347995765, 93.06929562288798, 95.92314482144022, 97.30200514749255, 100.30117871288859, 103.81270995442011, 109.89758484192602, 116.34876720814985, 123.89017747819523, 129.18672637515328, 129.27448751446568, 133.89403025842552, 138.96673300475322, 143.4434359406495, 145.53503571775903, 151.11992752295967, 161.77274701228262, 168.37833060608503, 172.65220538662422, 178.49559315547788, 184.98860617415437, 192.77759901009756, 204.73147346118384, 212.65664190547793, 222.78536445142748, 232.86075646846578, 238.92390046318346, 246.30108837038048, 254.1550211536378, 258.08230098239403, 261.13642321505966, 262.7320778035445, 260.07558238400594, 252.88428481826818, 250.39011261276536, 249.23151661613767, 247.72379039169698, 246.37638738145708, 245.77067318496438, 245.8389212141683, 246.01940224934302, 246.05136069945127, 246.20959341123378, NaN, NaN, 31.633496538360593, 32.14576489137414, 34.423194739606416, 34.49445968325767, 34.41345776010444, 36.39508684700803, 38.07852075762846, 42.117032359470365, 45.86090781178687, 46.81047493305338, 46.87517728679589, 49.36409751544387, 50.97093672642692, 54.04535162455079, 55.949186335540624, 56.38316309805032, 63.05940063633657, 68.70519471966954, 69.50985809817259, 74.3583250541715, 80.34110979725537, 81.21953702677874, 81.65176818673675, 84.72875687531172, 88.6841096577844, 88.24144280656915, 90.20995228684058, 93.06273877723365, 97.67746327149841, 101.1943467640754, 109.09741824847565, 122.51230733224156, 125.80957443485197, 124.27990344888366, 122.73217845520647, 146.9247873985465, 156.8220617990312, 154.17928029432022, 150.68813101618113, 154.02991423885928, 153.49118147767157, 156.7372340396173, 166.41747281868174, 173.9838279786091, 179.01714424847816, 185.039909829519, 190.2444968529108, 200.23691825185907, 208.8847612290544, 217.0711040863547, 223.53085723596183, 232.26832201078082, 238.54135085246185, 245.40852395635818, 251.73766839347078, 256.0937790868609, 259.99255354884133, 261.5355480557318, 262.86393170836004, 261.20131213535814, 254.31488424330536, 249.96318666173133, 246.6618198037461, 245.39067814800813, 245.53046316473635, 245.78372787912048, 245.67929117526378, 245.462230479666, NaN, NaN, 31.30306708569067, 31.557653455013174, 33.28404615540362, 37.14582706961721, 37.582467707570196, 38.312850941623964, 39.633789959350906, 42.3098081587331, 42.33896729995572, 42.80893700240308, 45.48713541490031, 47.100030632596635, 48.48844976701318, 49.62209949865679, 51.63728921741524, 53.58011811333307, 54.34460121412596, 54.51841561632744, 57.37629701015881, 61.22611830704897, 63.75324425047494, 66.17050598111683, 69.79582900690396, 76.83897040565051, 80.90915676994928, 83.87469610297539, 89.15256885543648, 91.67107469253234, 91.2268665507994, 94.08125211907114, 94.96719982689999, 98.26206365243969, 99.68624297724402, 103.41598209578797, 111.21674232149157, 123.41535823599321, 133.40719462019032, 138.36352338534667, 140.88288122525304, 152.21115017328378, 144.15830543345564, 144.49754732372497, 147.48357204816676, 147.531938283486, 148.3295852639212, 152.34992262075394, 162.8724291990563, 173.54451698853416, 178.46729952937486, 185.10457227037838, 190.33523183721812, 197.29705685905168, 204.85850700028075, 212.22067486905533, 220.9228288547547, 231.9122064581755, 238.84520004169806, 244.0023446866726, 252.38215874598308, 258.3011914142596, 262.4959635946603, 263.7834526643282, 262.8225436335475, 257.2915833132489, 253.1475802598832, 249.95485399583143, 246.72433693676692, 245.55019260430396, 245.1506020526774, 245.12055826189066, 245.0121348442013, 245.13675271929742, NaN, NaN, 34.091642897860744, 32.68974759098426, 32.17144816193593, 31.871160083593242, 33.41041414673115, 35.24524769888092, 36.19626755344318, 38.692755948391856, 42.441829897529225, 44.198458651083655, 44.70667817640187, 44.1851100678905, 44.25165266725061, 46.153490461027666, 48.79333099907243, 49.4506122243062, 51.13211027104463, 55.16238212346671, 59.12298238854097, 63.82093079799766, 66.05131219335944, 68.69121727088684, 68.80818997313692, 65.17258778111623, 74.85539096220279, 85.4130617567466, 86.17177347838279, 89.90671825337134, 93.30398352329254, 95.04743166531306, 96.78963516801952, 100.73787711735028, 105.80608017254865, 113.06693536913286, 120.65607617022037, 132.18020972545972, 141.7418992841218, 147.80596906875684, 149.5718874778277, 148.59774802724928, 145.76080924052383, 146.00999848245692, 154.4024381854866, 163.8266013517914, 171.9702674820596, 179.67372132810183, 188.73913695444517, 196.76515648215133, 203.34982746280863, 210.60218463561355, 217.86051993045663, 225.27546170171334, 233.31401890877802, 239.01222296592584, 245.34369286838034, 251.71198576197028, 257.4778436557865, 261.6005739031624, 264.9501502030558, 265.1650133228012, 264.70767081862857, 257.8678147200209, 252.34375840792262, 247.23222540922114, 245.2826075690957, 244.89696613421, 244.93372468874222, 245.03577578763972, 245.2096752821207, 245.3969381835468, NaN, NaN, 29.52778062349471, 29.155255822077525, 29.961654801882393, 32.86379379736933, 34.95428732909102, 36.23351759250955, 38.142826295689794, 40.48978852946877, 42.72682416692196, 44.30221258846779, 45.58227869802655, 47.19118797183184, 50.488584428245105, 54.11473909705038, 56.82724063643499, 56.855807192428365, 57.02901193580636, 56.797120547976554, 58.73541188970084, 61.33794871931113, 64.30464659412914, 66.50728300102145, 69.2495215986523, 76.18052661174909, 78.49237755634574, 78.04656084860841, 79.80944424494842, 81.78756076230614, 88.04812744037243, 96.84984979681832, 100.47911299872258, 102.4461511529296, 107.60536016415438, 114.4229363141963, 117.83005425045475, 118.92545828364585, 129.3759453303289, 138.06887517278085, 150.83036737349647, 150.84870069363637, 151.6295235331582, 150.5560679659862, 155.995745633917, 168.87202155006108, 175.5876510714079, 181.61933897326864, 188.63417234134056, 195.76476572015505, 204.3029510295694, 213.30232295843626, 220.52654858968995, 231.56915359260674, 240.13795535249466, 244.87127365849008, 248.6930371552714, 253.84834119162477, 258.57390445681557, 263.29208406656596, 265.1026744234319, 260.1069411032735, 252.866515743155, 249.79624164474762, 246.5195424196024, 243.9188899091521, 243.83369674029387, 244.10480302147855, 244.2676480894515, 244.33295554867357, NaN, NaN, 24.04104269468, 23.375328289860533, 24.549089864617187, 26.08788804438315, 31.74571661396798, 34.460866896238485, 36.29358333048944, 35.33271185958768, 39.14687007549257, 43.03870468508486, 44.06370314323697, 47.4389424489974, 48.53738247242224, 50.000011959433955, 55.13519912521351, 60.49518563784388, 62.84032477878024, 61.003389290802524, 63.12836892423001, 66.57117792164986, 66.93293233680333, 68.57741293098015, 68.90514270653806, 70.4304883195145, 76.36296826572634, 77.68167371380112, 79.87607156509809, 87.24482973126128, 84.82605630652581, 83.16606194043356, 83.8123316150441, 89.41716972675538, 98.76861418352098, 104.49563861022057, 107.67793625492008, 112.50994028880153, 117.4507612356293, 122.72931090324226, 128.02597204191238, 135.2823687471728, 137.80293500737068, 149.1689458499628, 152.6325647931886, 157.65378278233916, 169.51121975489835, 173.8314820400602, 177.205167643355, 180.76119514742211, 186.13648184179445, 194.58749231327417, 202.57925181042344, 211.89628402019693, 220.58750148543623, 229.34199784475746, 233.9216754203627, 241.47939135538834, 242.9785394412384, 246.17840050852294, 251.06768426048137, 253.01787722615134, 258.0840186691135, 262.44923832906636, 265.68239905511604, 266.03286225956543, 263.3893326428705, 255.30060394746522, 246.88426779611547, 245.08989961243944, 244.9838116760691, 245.1636278827729, 245.33259076003458, 245.43712371456203, NaN, NaN, 22.606287021387207, 22.30716079311692, 23.410536037779266, 25.248029469896544, 26.713845015277332, 29.79924838390367, 38.475739228655556, 43.39585658727401, 44.344547459885874, 43.52815367466364, 43.22744659520658, 45.936968285071515, 48.06001894284557, 50.477310337269415, 59.360554209960576, 61.487888457999944, 63.39541485819101, 63.69096852342558, 65.14662542805121, 67.12156498372364, 71.19170806225526, 73.16447662363551, 73.04632986985696, 77.76859287069472, 82.60097621830573, 84.68386693002705, 84.5718315344831, 85.00676559433441, 88.7434580021732, 92.48620003577427, 98.63771727457112, 107.98263346330613, 115.0124764474451, 111.37158735503722, 115.65146308898063, 120.6933436774424, 122.45710987212922, 129.9578532308517, 136.79082227804437, 139.64272289187124, 143.8708826569418, 148.9149138865549, 154.54702486137361, 167.97023699356873, 173.62824164823283, 177.3455823372911, 179.8049663310091, 184.03231095157474, 191.40889025915328, 202.84643936033495, 217.96811975221564, 227.28282194389172, 235.0045310272016, 241.73587334032544, 248.91256097526656, 251.9784908206181, 256.63969281194466, 259.80735419444574, 263.0267817557698, 264.80022286318075, 266.084087035704, 256.082844796045, 246.36691574846978, 245.310638121172, 245.4968386681793, 245.67469018914807, 245.85284914354, 245.92083023237885, 245.9922411055297, NaN, NaN, 26.811294012216162, 24.6712982707162, 24.29825867171886, 25.39573755292238, 26.273606403319366, 26.855998186131593, 27.365561122840745, 28.24175435146101, 29.194230792855453, 29.852422204174665, 31.169863871497267, 33.14918104202529, 35.495861727690915, 41.44494942899998, 46.72836516869536, 50.90934261881592, 55.68035582090848, 61.47611246011047, 66.0242985414617, 71.74892653768448, 74.79674467976056, 74.64088582947923, 75.23258106495318, 76.4685488688537, 78.80412142656783, 80.26146297876416, 82.8951637398042, 88.39188531185667, 90.8753563266732, 92.1087163752758, 94.95649832177827, 98.7519465668747, 99.62900401351153, 101.30865896972671, 107.83561068793404, 111.8624679837084, 120.50296029442707, 122.2074712266933, 123.97207380898101, 131.2309104387895, 134.87463856056965, 135.78713781701572, 142.42068926680696, 142.6449451321127, 150.49748590087282, 164.31262758156058, 168.7814588669351, 170.91080254666934, 176.5724586528739, 179.63128378787943, 187.4032647571007, 194.33261688824004, 205.29882367002122, 217.5333882461671, 227.87997245385398, 235.13732213038847, 241.2077326496029, 246.05466386523028, 250.03694930041758, 253.50158753180855, 259.00755386106005, 263.48384214687377, 267.04351373539373, 258.59493148643935, 249.302847498711, 248.25329769614035, 248.42100795862123, 248.70205915216846, 248.98530564540448, NaN, NaN, 27.200657319885043, 27.343267318846276, 28.444037763055505, 29.691696573360534, 30.86313933192209, 31.078257160147743, 31.513237304488158, 32.39142549665298, 32.90088460345552, 35.250587736823825, 33.922694923753774, 38.46970308069779, 42.069541005120456, 44.632618829582704, 49.98734299490977, 54.532540515303666, 58.85333312738315, 63.46989001258753, 67.35157294813762, 71.67529635351262, 74.97144127504018, 75.41140256882223, 76.73161438512516, 76.94830275801921, 81.34315219471452, 83.53934313652161, 85.28976948332873, 89.75734860091286, 92.97855969827295, 96.19131702014732, 99.9235262795584, 100.94802918100953, 105.27409614480126, 110.91192203533743, 117.81129844181179, 121.54154436795002, 127.10370719959528, 130.18403107791033, 131.73627893396898, 140.97786407979044, 140.93229781906092, 145.57972418545438, 149.76317313839385, 158.28954196460276, 166.27846636781064, 170.5383664113731, 174.6016812531428, 181.36102819438142, 191.48366791631312, 204.12963753880211, 217.08698120068, 224.9488033954651, 230.48969371036736, 237.2008548343354, 243.61774892162958, 249.08806307333174, 254.15139789336442, 259.7565128145834, 265.38780673676854, 268.3068191064602, 266.31221495066654, 257.033981175053, 251.24191481945692, 250.53016077668744, 250.69030058588797, 250.95522061813682, NaN, NaN, 28.166816564768933, 27.242416248218394, 27.384781233645853, 29.03488827082196, 31.6048124367256, 32.44903869275251, 32.40525806751114, 32.4387391738318, 33.754724517959836, 35.73699474288276, 36.577825428922054, 39.25393593417813, 42.92251325234153, 44.78913126687575, 47.28022042635302, 48.888857790034216, 50.60563985665374, 51.48566619259995, 51.77061646707234, 54.14965576193675, 59.61269994297885, 64.67105493810254, 64.9907855524122, 65.41665668224876, 68.16235438607269, 71.235089792654, 74.31080583092063, 76.39705869263899, 79.03411818598774, 82.43167329075996, 85.7274391617998, 91.3356427440668, 95.73288643354246, 98.25515876933837, 101.98310097600819, 105.9425246014232, 110.44991694251257, 113.41931291265298, 116.59811876653737, 126.50348079048965, 137.7273047920055, 149.39002549558998, 151.82922834257886, 153.29571853003503, 155.6585131581806, 158.34948284732815, 162.06429340133712, 166.764322427947, 172.24472861074366, 178.63374957893103, 186.70422924011334, 198.77109511652137, 208.6327428924667, 219.19539802665048, 227.52446506227514, 234.91500606473173, 240.62240219956948, 245.53324067726209, 250.437746341715, 252.14926815763278, 254.7868536175631, 260.1598882779236, 263.3415545269037, 266.3482972082337, 269.39936542024515, 266.10935395715853, 253.179534057684, 247.14185723309532, 246.87156713584417, 247.05107483470272, 247.2253285447948, 247.4203627305013, NaN, NaN, 26.029297520246608, 27.643303673675344, 30.658711790156858, 30.064556214386496, 31.6791556367576, 32.2617883082553, 31.887156493843325, 32.615177731608306, 34.226330859353084, 35.46977513365218, 40.605805420578506, 44.123286477684324, 48.672012140872276, 50.57606661400956, 53.50657739942463, 57.83469689805901, 60.254183077972435, 60.835590031071625, 63.25505254403302, 65.59311126758561, 68.67019645788511, 69.98338500621249, 71.84654053870781, 74.14028778398203, 75.89129530201757, 78.8560595776441, 81.93817478205229, 87.32507451681502, 93.04892066328013, 98.44423266834684, 105.48595805324751, 110.42045609211152, 109.32840562584215, 116.58906913199218, 127.26041677476678, 127.58968445118857, 130.2129534565793, 136.0363471246136, 137.23293771020076, 141.53165962472372, 145.72554894228168, 148.66620479358778, 158.36227680068845, 160.48494531771505, 163.05991518038303, 170.20990555833217, 180.93765273038767, 195.2773075490802, 203.11711800256128, 212.0358532490705, 223.7520101942114, 234.93471422606729, 241.07412595886296, 243.448374442016, 248.64549670706668, 253.50252467221668, 259.0069686442156, 263.26111359157915, 267.2441950370202, 269.8085492249421, 266.0162233774422, 250.9907465863002, 246.67028232912386, 245.9885730445822, 246.1250889080476, 246.23121574125034, 246.35658625526875, NaN, NaN, 20.795612400390294, 20.277199929713934, 21.010778358438806, 23.361018351216444, 27.110917542937848, 30.270976589989136, 33.647262638144554, 36.068101138543675, 37.683660005785576, 38.49431697843929, 39.22031058483314, 40.46067655313244, 42.3618022853571, 44.77972434686256, 49.400077815874894, 55.41711236248294, 60.32893548490772, 64.06272567010213, 69.71023864638865, 74.77314272678417, 78.4311477230549, 76.66172679754234, 77.53754998933039, 77.75522728842265, 81.4943261037143, 83.75754598264693, 89.54943760486401, 89.25141288644326, 86.09326909691137, 92.38810046244713, 94.5976652649522, 93.77884660942408, 96.99048442089665, 102.55451727200041, 107.52352725802115, 113.01404338622504, 116.59683894324642, 120.46244627832287, 125.80869255508046, 129.64957102562087, 130.6496130875836, 135.7181723744073, 140.6937601207572, 146.47877662900106, 157.9041046745606, 163.01558231138938, 170.1453691037641, 182.05019513036743, 194.1799841367396, 201.96364105702563, 214.12508350742547, 223.89438670777548, 230.23543061195517, 236.2442024068987, 242.17341369102445, 246.86623142246438, 253.67995064353548, 257.9624695684459, 261.59037788841033, 265.314253922781, 269.19794022900385, 261.61185997860764, 250.39153780245329, 247.72275494021662, 247.46927389210023, 246.93515022094172, 246.2625401682997, NaN, NaN, 22.129858566746044, 20.137864334495784, 19.3236536606433, 19.025567376934152, 20.197274071773915, 22.915835603460206, 25.853602281707687, 30.626600481106344, 35.474542986569624, 38.99891376113733, 38.55408347214241, 40.23594949578972, 41.70415345961495, 41.54840321435256, 42.56730525586557, 46.01214601553628, 50.04773087463636, 54.30426002003504, 56.27440617428115, 58.68579094698228, 64.84382769054096, 71.45157008266959, 75.33621271373335, 79.51264773077708, 82.73217241290388, 83.82818292725274, 85.87579684128919, 87.32720748462945, 88.71336308870424, 89.36803212100031, 91.77867963603568, 93.67485448927509, 97.26623994595911, 102.84320719501288, 107.31490561843808, 109.72301576548553, 111.91667441720486, 115.44094379028475, 116.18104822419497, 118.89651260061007, 125.76446442281951, 130.7582299706562, 137.35895078683578, 139.42538594628263, 137.54194205474195, 139.45697177186423, 142.26193835948848, 150.3923657516966, 159.86738058689116, 167.85770581406797, 176.47227788436203, 191.35313772624292, 197.32070368267134, 207.02245655426356, 224.61427326061497, 236.35937091868286, 242.85814469543635, 248.7730627945435, 252.59734993297397, 254.061748982578, 254.9095461292517, 259.381810153397, 264.4767680273438, 268.88946979089707, 261.4651843219024, 253.12014355502484, 251.3726362508528, 251.26180100655884, 250.08985370505258, 248.6347678016071, NaN, NaN, 30.04996504350589, 33.24802062063457, 35.011347035762476, 36.549748368586634, 38.19939843442909, 40.730393743690186, 42.708022583344224, 41.376917896395184, 36.85042104075266, 36.06811769779601, 46.97707393851234, 53.799384086527866, 55.76970993615655, 54.65913288001675, 52.23110552445721, 54.31466232085158, 56.07035895454713, 60.25422216701485, 63.883294558665646, 65.85147676208179, 67.9325551175176, 72.03334771192107, 75.91552031057616, 83.76096770383084, 86.7688095870977, 86.84069621192275, 88.52343783818536, 93.06184529289547, 94.22788656937192, 95.39517055360179, 97.71921464713841, 103.8689920579339, 107.96618461138172, 111.47986113319129, 114.78007690635451, 116.81724771444391, 120.76695619104754, 125.82833506188027, 129.12988653785018, 132.26950486156787, 138.59382739602603, 140.23165042971573, 141.00728199922594, 144.98128955141522, 144.14541601571165, 146.1648689523323, 154.86362878107565, 163.592555127705, 170.27120244442494, 181.76062902014075, 194.057907736912, 194.54764378789307, 198.94608197534427, 211.1220328863552, 222.81666017138753, 234.4384387400301, 244.073082249402, 249.1569218727992, 251.98901205625725, 260.0078947841916, 263.2148771001402, 262.1028496819656, 251.28563357947186, 248.60106124124914, 248.8829119260257, 249.19595529980302, 249.3628016362626, NaN, NaN, 18.405479005565173, 17.812830960442422, 20.09392502681497, 24.801917801547454, 28.40535877197004, 33.47849452330291, 37.29831656034196, 39.27829720485898, 42.579179162017624, 44.63214025595466, 45.735719225425655, 46.826319394515885, 49.093879097253115, 52.31813802092172, 53.47947237953325, 55.086860377373576, 56.91341669130542, 55.732845689989254, 57.854633349026315, 59.76364519461763, 63.688268300954306, 67.79313049947008, 67.4253375666248, 68.00335969986212, 68.43446332232303, 72.89799682745387, 81.32306173361816, 87.47090603081693, 93.40280441202171, 97.28306018998849, 99.62231734214707, 100.56122136863519, 100.18212628099802, 102.36939717768246, 103.82534090726622, 102.86500039763179, 105.72028990233231, 111.34805624155611, 116.60380364568339, 118.9339590104418, 123.5138733927173, 131.11888036188242, 138.0915186401125, 144.9123881577375, 144.27975042987856, 148.5930240876786, 152.47794111421413, 153.81925243991415, 159.07850081951588, 165.88754120783335, 177.5213566013794, 189.55568303096547, 199.4408357267474, 204.96131444594445, 218.30439410646113, 227.68361587411445, 237.44002302310665, 243.90704730561617, 250.94533473388847, 261.96186601502114, 263.70990824667837, 262.50885597496296, 260.61856440574917, 257.76153920998735, 250.97018201040677, 248.58062171750424, 248.67311201042273, 249.06379248665354, NaN, NaN, 18.73921161621657, 18.95659481587023, 19.173911575636723, 19.610113741409574, 21.001663196504634, 23.79230723378644, 25.113508695377522, 27.756525281832385, 30.25313777339186, 38.11456085589825, 43.47628613738679, 45.52522614393286, 47.64685141586379, 50.28688215067089, 53.074846225756666, 56.00539346867149, 58.78632573662992, 63.84304072508075, 68.09298049487471, 69.62243196409752, 71.04521736963922, 72.35305724627219, 75.98283732512044, 78.52059886896903, 84.23636493271553, 93.90182567038963, 95.98991953953384, 96.21341128798765, 97.4180723123415, 100.81195109805054, 104.53853038826855, 106.61629969454762, 110.79691411978384, 113.10711573587639, 113.98514920402305, 119.91855323664248, 119.6950388576246, 117.37994326010529, 117.93648221381146, 127.93051463076213, 135.32506803054486, 141.33858924722696, 140.74683765669803, 140.45349059316473, 142.23103344776777, 150.3244406932709, 154.30711790552806, 158.17737084977776, 164.73630245069222, 167.41460619995527, 173.4182112201724, 185.08922200404538, 199.505795073952, 205.61394677697618, 214.16404800150696, 222.93588179266558, 230.86266599401327, 240.09798933086952, 248.45337006622916, 255.7235632359781, 264.8791912319001, 267.4204508149433, 264.66997627846473, 260.4517174631636, 255.5050855866752, 252.2565654686133, 249.51251496107807, 247.3956618294958, 247.22862799035485, NaN, NaN, 21.976584958068347, 21.90543182406446, 22.051498905877676, 23.077279086234622, 22.561288399564386, 22.414987015623783, 23.51555359339053, 24.761550452772646, 27.036044620628566, 33.21309410315842, 36.07186246194962, 36.35238233567592, 41.930972730033886, 47.5858032663924, 49.93347894157051, 52.058205708900665, 53.95636716770342, 55.33886151744864, 58.337197738849795, 61.27261515980931, 64.42865447094717, 67.87453049311254, 70.9454055377012, 75.85326158249262, 82.16798254700807, 84.00161302415802, 85.45681826553943, 88.82677200801022, 90.21526459911794, 96.228873340226, 102.60978265230334, 108.84409913422176, 110.8099009990686, 111.89761874328705, 119.0869535979554, 126.62303444348339, 128.73035189360257, 127.029404290433, 125.85342548265022, 130.53090817297007, 138.7819285029222, 144.82887054475142, 142.96384864626197, 140.89632437296737, 144.41790616295762, 150.81107781918604, 154.79359461018316, 162.57721590730966, 167.92481430015516, 171.92885165988545, 176.35402201164405, 178.48454717543308, 184.56481316060788, 191.8481658926314, 204.84039594086516, 213.6470788058191, 223.95137275370894, 232.30786975946017, 237.89453755993233, 240.79609736035408, 242.9625047005039, 246.86039431263882, 256.52599602700735, 263.76833436634365, 264.38161854537174, 264.6336340338785, 262.421020564265, 252.36326011941725, 247.31670935799968, 247.16149488911677, NaN, NaN, 21.089024877548, 20.31517830202727, 20.7573150655932, 21.565995375272685, 22.077363227400525, 22.917536318475772, 24.09088675215128, 24.67387239555359, 25.22039176739642, 26.13566145999547, 27.234197256677522, 27.961636774780853, 28.144129643225757, 30.458517513760064, 34.09651744270686, 36.81459243197764, 38.60989516562365, 41.06812440742355, 43.11398293993416, 46.99979488008568, 56.75975104247655, 66.76819543594083, 73.48114346972915, 74.89211769498452, 73.57386520617214, 73.35073049829398, 75.21387548028855, 76.08083640391362, 78.28288318008164, 81.5724555720848, 84.53087200989283, 87.26611555560987, 90.11478212659898, 93.0876743720482, 97.9257019607643, 102.20050640594422, 108.025546023324, 110.65751919254066, 112.95982452075059, 122.63294248883284, 128.55837070086216, 137.90331561824257, 141.84305191499195, 147.23002779665973, 152.37923345775656, 156.7538228369959, 161.39578127245008, 162.41100314188412, 164.96612060259744, 172.91926381976324, 176.0365931146898, 183.4790314596469, 192.1501746034203, 198.07024952691094, 207.51790571402105, 217.02621683737698, 226.4323017364563, 235.78956305692253, 241.4550859690642, 245.76675000885513, 253.63734981768437, 258.2594257932186, 263.98805693953943, 265.92603652380734, 267.04390469779867, 263.9937773950891, 251.84477848304365, 248.1465088777121, 247.99930458991426, NaN, NaN, 19.607965574415985, 19.345869393509787, 19.56260525035304, 20.442467872365583, 21.246872539524745, 22.753752803125007, 24.331211465335837, 25.022602617450673, 26.122011422872813, 27.51504342055203, 29.165223603591095, 30.407496214905414, 32.05669583631533, 33.631267470818166, 34.76375308538763, 36.00458783683435, 37.69006292522329, 40.51822651255123, 43.30508378482311, 45.616752110959766, 47.406921836083725, 49.458465681222485, 52.530709066869, 55.38479042448836, 57.288104459885, 59.036389735121716, 62.11327024713147, 66.73273412715199, 72.8928309760104, 78.31874321608221, 79.78892154161144, 80.28598914555755, 82.54548216291761, 85.69685020506155, 82.1820603684846, 83.56072953704624, 87.65457436971921, 94.67751871612928, 98.19598152520231, 107.20664980054408, 113.00231106042108, 118.70059339886656, 113.41668922802157, 113.62137849133018, 123.0008102291143, 128.67853993584015, 125.5828412501042, 126.71365673438308, 131.33942739543113, 149.80358548511427, 171.4450866443104, 185.9629517603333, 199.6699650295005, 212.89278658266954, 225.4483811919059, 231.29482405606032, 239.3975518175794, 246.5840119779616, 253.36964313788982, 262.3084411688517, 266.29606517935906, 263.7126871497768, 254.7573817797769, 252.56569851908304, NaN, NaN, 38.46833127241159, 38.130720914312626, 38.41601679921526, 38.91843091840148, 40.12460614827517, 42.9507025241002, 44.85634618113227, 47.64618640023747, 48.99464346638663, 50.67831279398426, 52.68942997817896, 53.73839390183618, 54.4192676673658, 55.62168977746144, 58.780052763347676, 61.379236971716296, 63.75575717500899, 65.5761991556367, 67.99530300852663, 71.88447249273977, 74.99528618980214, 80.28292800536373, 89.09064217819399, 91.06908261665161, 90.39903122082481, 90.82840268315924, 92.8044652437819, 94.78477248805763, 99.64541441429934, 106.05152370411486, 110.26170021053777, 114.90433422795434, 119.78041039493434, 129.4847302220008, 138.99264760371872, 142.9685045811662, 143.20946070740854, 151.4882395484481, 176.95896703895014, 194.84843248310392, 202.47419479947138, 211.20530110032718, 231.26369098469732, 241.51340805258317, 244.43837197499744, 248.279959793059, 250.72379045197354, 254.60750586996542, 259.37413741101545, 264.8150168819645, 265.07392181120963, NaN, NaN, 46.145817372602295, 46.291378184545536, 48.20221139515465, 51.51340559889383, 54.300957230090724, 56.868100657239104, 58.54785440688222, 59.93197394655129, 61.17137092134487, 63.295402990272976, 65.33923210677634, 69.01756707797796, 74.45287271830554, 82.09781090328745, 88.32846696488664, 89.57584231815461, 90.2481735995475, 94.67736871107967, 98.6346467855901, 99.79908129588725, 103.1319232567384, 106.37500193322751, 105.47859838190824, 107.85274351403373, 110.81606739119216, 113.14460782951238, 115.47870642795439, 115.25153645189835, 130.907712487743, 165.46943363886692, 188.14385987015152, 199.07257026706353, 206.79123856444784, 209.44656538084084, 220.6566969772383, 231.4885769241386, 241.83270443637034, 248.83574833733832, 252.77362425527218, 256.38774351811986, 263.73490154745656, 262.816315650571, NaN, NaN, 67.92938373194796, 68.07492066792874, 71.69688527999631, 78.24991827142142, 81.47476400390804, 82.99490973353876, 83.55916248728286, 84.57723144792595, 87.3709158521027, 92.76129699805864, 96.20443320700306, 97.80837178422443, 98.24773754400663, 101.0950987641126, 104.10014454925711, 105.65788984614392, 103.87150027778311, 105.12058545221043, 108.12122188588488, 111.54731829212412, 134.99460215824874, 140.5202145538731, 142.89142410845966, 157.82099675958128, 187.7034251283239, 198.54151176793272, 206.85602629425745, 216.59848714910567, 229.54652937646944, 240.68147058305706, 246.00261053007299, 250.56522589708953, 256.39661935045126, 262.39787735700503, 263.05869318459713, 262.4445855613766, NaN, NaN, 87.42738919685426, 93.34550058020139, 96.29981558483755, 100.34965349630163, 100.70082549076537, 100.68314104695166, 101.018178549026, 100.98620893802962, 101.70292223356223, 102.78992375285185, 107.55532274786854, 114.89159929991376, 126.6813056913662, 134.57689273238103, 138.29241439542616, 181.7536303621422, 200.92032156251315, 206.0753869387601, 211.28622036686454, 224.168562254687, 238.07848124137553, 246.60359780540747, 252.1792026915027, 260.2448909389708, 262.9267613275018, 264.20533585276684, 263.37060218380014, NaN, NaN, 95.22858864452033, 96.22472104984669, 96.87910232704603, 98.1936934656713, 100.1625646157845, 101.12913523274861, 101.09965519893633, 101.73955197641189, 101.39493202263121, 102.36217132520257, 109.29941271812143, 125.17373992789888, 138.13525276248697, 134.35248209717116, 174.1749005098026, 199.39246101449376, 207.01508737029516, 212.6821929775296, 222.19106329354133, 240.17756196197868, 251.02475719932664, 257.0101580076096, 262.78603588306026, 262.43806468899106, 263.39415600267347, NaN, NaN, 96.66095641411879, 97.02269986632629, 97.74324876093314, 98.45773525075235, 99.18468183961234, 99.52681262306946, 100.96476223829431, 101.66675950934025, 101.28357601625426, 101.27120785936813, 103.09236170645367, 107.48213170274711, 131.41232462991587, 139.6617503489869, 143.43508570794813, 188.02821804738022, 201.263821828877, 212.02941323407708, 221.79420316063306, 234.38134034273386, 247.50727993529063, 261.3602536637092, 263.9010123777079, 263.06634865795, NaN, NaN, 94.45637183189292, 96.22724535507753, 97.09131614709158, 97.65636951401721, 98.22046895354592, 98.78640192232638, 99.35081155387346, 99.32900660093115, 100.77102718108117, 101.62971013915984, 101.62106209970071, 101.90268046950501, 116.33319955060297, 136.9595482917022, 141.84562841330964, 141.60406926322125, 178.77519746851567, 203.2826818720777, 215.85416630897018, 223.30962500437568, 229.90825883824488, 241.60085742795826, 257.59389073202294, 263.95444866319565, 263.3967503884105, 263.7987711968497, NaN, NaN, 97.85479261954295, 98.17470702563861, 98.1553224683436, 98.80712826652707, 100.12505317250478, 101.09083759258522, 100.72847968504502, 101.02732187456381, 101.3334649706278, 103.97271225469535, 123.18846526359336, 143.80785601867754, 146.53646149148662, 134.98990236990633, 154.52424806585566, 194.36503167846558, 215.49362711214584, 230.7180319779125, 244.24791776477736, 260.5898303241615, 264.4966389082596, 265.0426406908811, 265.16710627445804, NaN, NaN, 98.39931012619607, 98.64825852803577, 98.88700229716855, 99.65292580436525, 100.41276043870337, 101.68335318111039, 103.20763525906368, 104.98261203480435, 120.68190918630093, 139.55600264477897, 154.27947539390303, 154.53227770894154, 141.44534219712065, 136.8059360598297, 152.49447793332726, 184.9344792052731, 202.22571090461588, 209.25080513984864, 220.60092957249583, 233.5345468281624, 244.01075653246383, 259.7072022454674, 264.0583354972965, 264.4797936693844, NaN, NaN, 96.47579905436598, 96.91918756448334, 98.46611191256538, 99.10616729516299, 99.52568699516783, 100.16487279246263, 101.0385588433879, 101.89563592187764, 102.31673172341624, 103.40100279428962, 109.32480122809892, 116.55505272301694, 133.15811911155154, 152.48020209468893, 143.9786107295911, 134.03537756814478, 143.51248909093408, 162.2334967784695, 187.3961707456123, 201.34966882437692, 210.7478937346067, 227.36459888754254, 240.0460017715127, 255.61320729999932, 264.6381623483835, 265.2587957795966, 265.658642611999, NaN, NaN, 95.69822245045512, 95.39490852453825, 95.67261438911362, 96.23715486893175, 97.10866210442448, 98.88804116782842, 100.34448275699683, 101.20092408744249, 102.50544765427638, 107.64117476092731, 113.05189484224377, 116.39596530993123, 121.65395897081126, 130.29632960274006, 141.57668237853812, 152.64019128075273, 154.3392570400083, 140.43391026871015, 138.35058083337572, 151.4130718615107, 175.09823464054068, 189.79722442159775, 203.30607576033768, 223.336599530575, 247.51487757452324, 263.6898633914542, 265.420539606153, NaN, NaN, 99.08431171404037, 99.51601875339301, 100.16373747256642, 101.46706069286016, 102.31305659184096, 103.1600389092891, 106.20864500558697, 116.30421334688535, 129.51422427304422, 133.2087860384981, 143.47463121700238, 153.72167343434703, 147.35721510168216, 137.22403915369884, 141.16758971134803, 150.63291398045394, 174.00003876690656, 197.59356361201444, 214.21372562478228, 235.30256892760755, 259.58354801679906, 266.4216314104956, NaN, NaN, 97.40999896443742, 98.32129885356707, 100.37710790177668, 100.93752601654111, 100.90841757151912, 103.22652539177064, 112.88381489390399, 114.02770602856538, 116.3563565439355, 119.88602426843781, 126.91342735306, 138.37409629533852, 143.09864044154577, 149.35642762592124, 150.3034224703675, 137.7347239557309, 137.72594810683762, 150.98379113251903, 183.9566916789595, 202.55274032210664, 218.3338582098963, 231.91244760215477, 241.46850948837525, 246.7918147699203, 257.45696531772, 266.53723313269126, 267.9258379807606, NaN, NaN, 98.92073963538914, 98.2393026496131, 100.67859179932925, 108.16395519485022, 108.58412328850376, 110.0971986792147, 110.94146252245561, 112.02609464691497, 114.41914930544468, 136.48127955270363, 130.89732011085044, 124.78188471921482, 131.37341224271077, 144.62424317590202, 162.2701316748287, 188.94557575141408, 204.88338715932633, 214.1037211977879, 231.9141590429724, 246.46330397486886, 257.4749264406608, 266.548054567549, NaN, NaN, 86.98932908970549, 87.59806031660786, 97.10213982534171, 104.74184280355131, 108.25552964043162, 108.51886038766814, 108.78561122759619, 111.13037876356327, 110.82337486127376, 112.28133302779949, 121.12577010460343, 112.39684057533171, 111.80758775628279, 117.10267840471985, 130.35950174298011, 153.91422328798456, 188.92535693674935, 205.5010796385965, 220.8504232400562, 236.93135756036133, 250.67612441792855, 262.54327996003843, 266.96269587045236, NaN, NaN, 102.08019959914704, 104.40888710137828, 105.9445124992238, 106.17605119346294, 106.92715365683745, 108.96466301571192, 110.994583258293, 111.76988675810689, 109.95408025566962, 117.17047914622158, 110.5515031543091, 112.1395026151006, 125.29418172119307, 140.2220267946573, 149.71609535722203, 166.42657798332232, 194.74921160690474, 207.45738118085126, 221.4204905304057, 238.83479564186385, 257.527090153706, 265.27012436996824, NaN, NaN, 104.9709489675847, 105.25619284049247, 107.03126889480743, 110.8253859039873, 114.03034968983933, 112.56897311589528, 111.09217547033825, 110.7649911674219, 112.50583421313797, 111.37016383352959, 107.86042156568682, 112.00132911742024, 118.16201591977591, 128.45392717657685, 156.41221309395297, 191.15968032204867, 206.22262965261206, 213.6944013867365, 227.3437400216673, 244.2538833578523, 259.9028104508105, 265.70206431502555, NaN, NaN, 105.0365653241239, 106.48988244810454, 106.51090734798863, 108.56596756714488, 110.61931506500831, 112.07822939304347, 111.18612268734705, 110.56290656420212, 109.68815457112989, 107.07481596607812, 110.6135240921092, 116.77853359781759, 141.23904743633972, 175.35153741177996, 199.8529610446205, 212.9376216333435, 229.10662586513715, 250.78719791949368, 263.29818193043326, 266.91751812419625, 267.2705830500124, 267.36722084798436, NaN, NaN, 98.56442322467204, 103.75241908371808, 106.60482903428225, 109.44146356279214, 111.76645429803685, 111.75915225771914, 110.95528043511041, 109.13080000772806, 107.82611853452623, 106.81587884866117, 109.90762834462842, 122.82412696286485, 140.5865811858545, 169.67616922151802, 198.29734843012594, 205.7782071545303, 215.7664958241476, 229.85889558470225, 248.99578698582098, 263.18510670924206, 266.21428199547586, NaN, NaN, 107.74446417446538, 107.13582167698155, 106.26392116909331, 108.33854917223938, 110.4058698672543, 112.77534201513863, 110.98677554056937, 108.61139266697884, 107.4134607722439, 108.58892931367208, 126.0659758642154, 161.6943777555289, 193.80567367217134, 207.99146989490063, 217.31918733931877, 229.13701597582863, 240.34228618554582, 251.6636545221007, 262.86077648980404, 267.0806960370882, 267.7001416065045, NaN, NaN, 98.55706557589085, 100.88503225883798, 103.72304681033056, 105.79475260093574, 108.89102460489721, 110.70598576950992, 112.76263671011283, 110.93259432845491, 108.59183800893238, 107.0298878356077, 116.62342272703366, 140.87605718450686, 170.46946832330192, 200.7454126920669, 218.0487961189567, 230.457516206145, 238.53803166059492, 248.0304722437297, 259.5018236960558, 265.2952964486409, NaN, NaN, 98.41355540609358, 102.2554280806513, 104.29858769704802, 106.08746772420515, 109.04146380878132, 109.9246747977745, 111.40200577068732, 110.81167600782996, 108.73619830691062, 108.41463813270728, 109.57587961785333, 116.68921146853143, 129.93407843465505, 146.41773756933475, 182.05006395717095, 206.0664809098741, 223.9278122342906, 238.93541514801564, 251.23108229827255, 264.18055112476304, 268.06005826796235, 268.28134933070527, NaN, NaN, 103.34222725629493, 104.14167125683664, 108.29394322113463, 110.3757540617775, 111.67359126962643, 111.64404802705138, 110.33919521785438, 110.34166747760956, 117.82023636794943, 123.75032024701058, 146.4252411271907, 177.61222760728472, 196.13181635336744, 202.05157516965096, 210.47730920733196, 223.556620564834, 237.65918380013179, 248.08985604750964, 257.9921985457231, 264.2453817428711, NaN, NaN, 101.61786327742476, 103.5922537704335, 104.56425039798236, 103.88262035968589, 103.54110921538359, 107.87908801666383, 109.85344521208998, 111.52946206146152, 111.84774084576316, 111.1640714002827, 110.85330034761468, 123.13722181918438, 160.61093015605303, 193.38992987874684, 204.78241343027992, 211.18860098136298, 221.05828184867968, 237.3176517643552, 252.08623285877079, 263.13321282171313, 268.3832586019543, NaN, NaN, 102.3766330314314, 101.70371784649846, 102.02438227115324, 103.99940687992586, 105.96978983383053, 108.29088621841125, 111.25548441264914, 111.8920325108821, 111.8672726853011, 111.21713825702193, 112.19129790516745, 111.84594941054144, 110.88628087948112, 120.49159767562105, 160.58627123716684, 200.16438886579476, 223.0120121091431, 246.42642322206163, 261.84967249835694, NaN, NaN, 103.11818907751618, 102.522355454739, 102.81195494230853, 104.55347490274801, 106.31130476683191, 107.46952981946248, 110.11081748033509, 110.96492930893731, 110.93171448555512, 110.62622682932809, 110.63712006894119, 110.65407570587732, 114.48734526253615, 147.5023923142958, 174.84552340617657, 206.5236799432191, 235.09374786251212, 258.87306561589304, 266.71520675581996, NaN, NaN, 102.93697362863918, 104.59490664303057, 105.23635561740724, 106.55434519483381, 109.18262680404591, 110.48247727065228, 111.1129122376716, 111.0784124213492, 110.07430504912207, 109.41803911956275, 107.76953811754368, 104.13645595462152, 107.12203281411627, 134.29887421337025, 151.17524667152836, 180.0095242969797, 219.29787756169563, 247.91475750490258, 260.8031427437403, NaN, NaN, 103.39287552685362, 103.38028007880743, 102.26652287698629, 105.19754264690309, 108.13497455477541, 108.4852878076266, 110.30244334070606, 111.00614964724629, 110.60864234440709, 110.21793721235802, 109.49276810743017, 106.55769390583517, 105.11654087915274, 117.62432862289319, 144.14646892295252, 189.45052444627834, 221.58925907935895, 248.6361607077822, 262.6905349909218, 267.2342875625804, NaN, NaN, 102.05954397542865, 103.2468448205422, 105.59664101918321, 106.17867773231046, 107.93995466059195, 109.97983160540616, 110.8283300260711, 110.79969664543138, 110.76716366732315, 110.15048519590285, 110.12717269417456, 108.96407934329952, 106.94236465857283, 115.81670295923833, 149.6479934529277, 184.34341031460465, 206.54650188742468, 231.7128971632196, 249.56945129064025, NaN, NaN, 99.8535302543299, 99.02389495908193, 99.82358288760135, 102.64945274981656, 105.05031049209032, 106.2460238837984, 108.66988296305017, 110.66313312910862, 110.64003290509415, 111.02427221735024, 109.00338276569003, 110.63440807711022, 122.00337293418849, 169.6442803610893, 199.3312166949068, 232.47819131387345, 254.45377040628765, 261.91194413240635, NaN, NaN, 100.9992640901219, 101.32084975655658, 102.62955133219937, 105.92500874197304, 105.91745503497155, 107.23643547728643, 110.1951077825169, 110.82696007207996, 110.47063740680572, 108.49411372000561, 109.49645432119343, 112.80302364556522, 144.87432594241258, 185.84739187838107, 204.20255647341278, 215.29664310641692, 244.1521319279936, 258.64315506405757, NaN, NaN, 106.29773222487131, 105.94468612644945, 107.07704225985351, 110.0202311457536, 108.58780577644626, 112.63423723824403, 141.728421589364, 186.61513452502595, 206.69516808860593, 215.61475480514352, 223.34403670461847, 224.33739418992798, 224.63649274650894, 226.0618153232935, 230.81260879253327, 237.09211397777142, 250.55830896771235, 259.1115808418514, NaN, NaN, 105.73657989972429, 106.9777078483005, 108.98996440973414, 108.98457713648985, 108.97976381855325, 113.00435618879844, 126.7462658111166, 176.48506769682783, 193.06821142932625, 200.85058360576213, 207.77674104025868, 212.6247769868738, 214.586806728355, 217.42193021175794, 232.56968428464174, 250.0648162823371, 255.33913373343688, NaN, NaN, 108.29817176643125, 108.74142853870978, 108.29704883529011, 107.40500596994696, 111.34788703309688, 121.02345510640713, 130.49433353826117, 157.6359231893632, 185.4494245071219, 194.7535024684819, 204.83544629950842, 210.5827406528242, 212.51231354595592, 213.80440047619797, 215.344923389135, 217.75203822365134, 221.50655649628203, 241.14485214336716, 254.94256522494294, NaN, NaN, 107.76996595562643, 108.21699152769168, 107.77060867230603, 107.30523803881991, 129.09282636092732, 156.16839413680404, 176.91437789358872, 188.17159975589345, 195.282585012183, 203.06527844643054, 211.53262345195395, 220.59733674219564, 224.13386969861043, 231.72152887772674, 248.423883750041, 254.90962326512627, NaN, NaN, 107.30226977309458, 107.2923707708845, 107.52947668790212, 108.03337576719748, 107.76703206315477, 109.54864059569154, 121.59837585141511, 151.62128612557834, 175.50951316828642, 184.80722057918317, 191.01832962971858, 195.96176172969186, 206.94730630138957, 221.9594095919523, 228.6707171148887, 236.46389713154576, 246.07251974142022, 254.73104256402888, 259.67755758287285, NaN, NaN, 110.21819034756685, 109.43123967946893, 108.64865055143073, 108.41757917022228, 114.83890200795715, 145.9263486675389, 173.7279471122655, 185.04068848991378, 190.45780846963672, 194.05031911517344, 200.87315135451257, 214.910183400992, 225.51244383369064, 229.88529188530038, 232.19621280071647, 236.60851951847155, 255.97523587380135, 262.6720085888284, 264.2208348207141, NaN, NaN, 112.24464714882473, 110.6837046246181, 110.91409548079422, 113.46744711992457, 125.01827372628287, 157.43643700300703, 179.63466758774325, 190.76295661129538, 196.1561900503876, 199.253950830635, 210.2189041584226, 220.3285371876261, 225.45083553038185, 230.87704594492897, 250.3838319764423, 261.3180669682215, NaN, NaN, 111.73625714028185, 110.79885011361603, 110.77064964598345, 110.92204174752304, 113.64390775194998, 131.05713471817128, 149.40878182563802, 168.7289821230551, 183.68894320761868, 192.3784433245518, 197.90829049067364, 201.7845343000031, 207.9233197712575, 217.93039480269567, 231.8324087597706, 251.2642688234355, 258.62975129634594, 260.44657304500345, 260.8074247332827, NaN, NaN, 111.87907189750331, 111.12316442408144, 111.28206998482125, 111.43341296538178, 112.68828464058576, 119.08138288807068, 139.98549308054012, 162.0171407230519, 174.91937459792348, 185.60563830357708, 192.4368014220633, 202.75118344150084, 211.93366889815795, 219.31607846608466, 235.07498192983417, 254.15218974620413, 258.5516466504439, 259.08879007181025, NaN, NaN, 113.9419213769469, 111.72012331333494, 111.50997791489998, 111.11377381069063, 111.09243193893113, 118.60216529558109, 133.98124057636844, 154.90733348202696, 168.29274073786073, 175.28874905961987, 183.407158248815, 192.74242357407854, 203.87398389175553, 211.42114053549983, 220.27384671623523, 239.53988624264744, 255.69391670559034, NaN, NaN, 110.55098592499232, 109.87052138881316, 109.62459873884357, 109.80998808572018, 110.00422169555095, 118.59274179683287, 141.70786202954753, 168.56792929381734, 179.87983699891288, 189.4798684208887, 200.82020780652203, 210.12477524745591, 224.97858492466037, 247.0013701851937, 258.20823876918814, 260.8402551577359, 261.27278701413, NaN, NaN, 110.81578978031342, 110.2803690641568, 110.25360641742313, 110.21284520736451, 110.42930813369725, 110.40421701157297, 118.35834629363461, 148.642407797374, 173.59487504193228, 185.59567953223308, 197.01151360547448, 211.80388733232454, 227.02543024996586, 250.50065284686318, 260.75205319158476, 262.53873148684795, 263.03984497157273, NaN, NaN, 111.31508283103564, 110.74333842283497, 110.71985792262159, 110.87149702202314, 111.94950081572475, 117.26065884515425, 137.05775821603623, 157.21729780406298, 173.56745423304838, 182.45987978941548, 190.0730610230752, 196.91726300946883, 211.78349962431173, 230.99010080027637, 250.29291754493613, 258.805367149845, NaN, NaN, 111.10984874014335, 110.57314707820082, 110.5448988778749, 110.50523974347858, 110.21590269559718, 110.72934066740854, 122.78060084330006, 138.68952184416878, 170.52743508207004, 181.41948294881803, 185.07549917004476, 207.16163877128105, 237.1835367512835, 256.09788541836105, 261.3253246168787, 262.3568753050481, NaN, NaN, 111.38901419541483, 110.63227151322683, 110.60519741762616, 110.57336054822018, 109.8229697565139, 108.71501596761415, 107.9701641694272, 120.8074670308874, 162.94695211322923, 177.9983511340441, 183.5854777293405, 198.52636629592868, 233.30470243969103, 251.8329378421686, 258.66525007009915, NaN, NaN, 111.31010561431852, 110.95835414105547, 110.93274315695619, 110.8969980265645, 111.87036104538689, 110.8627610510979, 107.5609686980473, 124.69554281587678, 165.60174713530074, 183.13956297668508, 187.24780429342894, 214.6628875981619, 244.6455296885095, NaN, NaN, 112.6201560743015, 111.13526074531228, 110.81979476972667, 110.78584349389018, 110.74778325579685, 110.41604780556635, 107.20504842187388, 108.6662067056555, 138.57231470533796, 173.71720126049956, 180.00007638743335, 183.33546712881375, 197.55839713803002, 219.53795822932426, 242.19521912196677, 256.7346303905283, 259.39285696507903, NaN, NaN, 111.25081482713554, 110.9761762050852, 110.95145492694934, 110.91516470891635, 109.85516040994764, 109.33163427881126, 112.43012879866109, 121.64298438350755, 134.4344308065101, 149.80667716966275, 177.02721540317964, 182.21306240337702, 182.89547231374058, 191.65346371854866, 219.79105547907267, 249.42105943394475, 256.91462027650795, NaN, NaN, 111.87856532682811, 111.19750640137488, 110.83809388675772, 110.47417683468052, 109.77750967002468, 109.74104635677058, 109.05935253727735, 117.00289359028179, 145.68166511093494, 176.36894878789192, 177.8706831542023, 188.8729248377757, 207.85312568722608, 247.0659774455222, NaN, NaN, 112.16763723765193, 111.33705453273905, 110.90335618078586, 110.46027630875162, 109.61280038661418, 109.20718942973674, 124.94148452689767, 171.7206621009787, 180.6785392318588, 184.07813523418994, 201.12750048997694, 218.20499055085568, 248.64637390211186, 258.4446535388996, 259.6587889058176, NaN, NaN, 112.2147596222993, 111.60444970141354, 111.28035997717667, 110.65258453131717, 109.45660525385871, 112.98969158481816, 138.47272954139407, 174.53249341726675, 185.71800495938996, 184.42067749223597, 196.0446123857805, 214.32929400304184, 235.65193510711322, 252.15130721736696, 258.72097810231196, 259.584571509046, NaN, NaN, 110.92369387781777, 110.17039100189496, 110.13790110537238, 109.73307389317404, 109.33920745409543, 109.32392853546551, 124.71766829361066, 170.88877420763734, 185.98593955301388, 187.13350923501162, 192.53341764516378, 215.11890006130182, 239.9002781078894, 251.5713967821157, NaN, NaN, 113.86742849907088, 110.50698969816021, 109.96516364735847, 109.93033260349621, 110.14965083207179, 109.6060516798001, 113.96769988103821, 141.64075195180905, 170.6206177267064, 185.62948696240446, 190.00533270171988, 220.12312348574335, 245.7191695879626, 254.91883327484817, 260.4705844833953, 261.49544284782877, NaN, NaN, 111.18450144340795, 110.39269527969067, 110.36134862723598, 110.32058254948834, 110.79529487962088, 117.9802775933833, 149.26188938732122, 178.29736334087013, 186.88532099683357, 192.48903556983888, 217.3990030101453, 248.52397064975648, 259.9681652207744, 261.3051540696542, NaN, NaN, 111.64708970105728, 110.96343669867443, 110.93616019729798, 111.22585303088566, 111.18677743042612, 111.48247369624353, 115.76945706607465, 156.37501346430972, 184.7827066469162, 189.5803264613878, 198.65889114542395, 221.67652139968257, 245.31583496006502, NaN, NaN, 117.04875257346575, 112.07457413520704, 111.38999050174915, 111.68720018814552, 111.65682102298176, 111.29599278427571, 111.26912365727655, 112.57716168103154, 152.5147228577836, 184.55793575764883, 189.91049597281634, 192.7463647834735, 210.48309950309, 240.4004330445124, 259.46541927029716, 261.49018760100876, 261.8249916683841, NaN, NaN, 113.18172414587464, 111.51092121353105, 111.4880595942882, 111.45747245160074, 111.42381221625922, 111.39961424086526, 145.74426114950876, 183.74795764644497, 189.48162735985673, 201.6483890276518, 233.89904719277422, 252.99628179024444, 259.670309231493, 260.98760860209353, 260.9880138863595, NaN, NaN, 113.92936482815367, 112.91461532000879, 111.89388160506869, 111.20303541761126, 111.16806758893559, 111.48292396282652, 149.81447405620915, 185.50347436042782, 190.61264973783202, 212.73624028937624, 241.99681437799205, 251.05893782181144, 256.0597432455592, NaN, NaN, 124.59187252670522, 113.99766881750347, 112.20667622652417, 111.72495566002081, 111.68076087480905, 121.35506675005962, 172.8863341032416, 188.8044168964081, 198.7601874449596, 230.72627497038252, 247.24116565636504, 253.8768728482742, 256.5376962066589, 257.43092436589876, NaN, NaN, 113.80518972600665, 112.57054641233975, 112.54415343713198, 112.50558708840445, 112.47436697243981, 130.6141781936844, 177.8633838246941, 189.27247608400873, 197.16134922682596, 216.6679220071792, 233.01423018984391, 248.51635443651836, 252.98648044035636, 253.4383304956621, 253.8660791604176, NaN, NaN, 114.53037118026948, 113.1856020098415, 113.15749445690048, 113.11349341043721, 122.78027711386505, 174.3387353777673, 188.94058470389672, 195.3149322043104, 212.20984762756135, 226.38721011189344, 243.7901491455219, 251.36023417314058, 252.30913415475075, NaN, NaN, 114.66067387379954, 113.4257538320482, 113.39513619559581, 113.35396077765785, 117.36998948703611, 165.79681827920814, 188.09107021332454, 192.68602219848066, 209.05309387864224, 229.3361974833366, 246.50446519615394, 254.27846185730687, 255.92029300755198, NaN, NaN, 114.94520773688684, 114.11687790287112, 114.09253385510645, 114.05221329527792, 114.41857451338696, 127.70763123211454, 175.77412682571284, 189.17110703713175, 194.62503386889048, 210.9561124287344, 229.65315687492313, 247.14377511803713, 255.24675319414195, 256.93286717680417, 257.78635875006495, NaN, NaN, 116.11350862524712, 115.10043940103694, 115.0705321456702, 115.0306140527306, 139.10899601356172, 179.77127954754246, 190.7894535597383, 203.29052752832317, 217.88781949654364, 239.5434834582646, 253.1745282701718, NaN, NaN, 116.36353703138923, 115.35107263840422, 115.32351077579342, 116.28788393942108, 145.33006533332033, 182.7022308813827, 191.78983232522626, 205.24781572512893, 218.83728865297292, 239.14799415854083, 251.47605576378703, 258.22913139906257, 259.87305386561144, NaN, NaN, 119.1928729893667, 117.15295594126974, 116.31736055932865, 129.63849927736362, 178.96455305312867, 192.9045771816183, 206.8468736016321, 219.78937178504643, 229.87997830382463, 242.51964956525353, 250.30511598756615, 254.8778202428172, 257.3250730893963, NaN, NaN, 119.64590942538857, 118.15984942362039, 120.19673649689413, 119.8802837962744, 151.62168649555176, 185.7558313113489, 191.7455062704652, 201.95029781061308, 215.24886864357595, 223.7733405567214, 239.49499263734614, 246.8891334006322, 248.99012331404842, 252.96386641454527, 256.8305170093284, NaN, NaN, 123.23535364103924, 118.81208511580715, 119.15393459389846, 162.13266363826352, 185.73769305086714, 190.61210625256834, 208.0330944036761, 220.50905490119524, 238.6137525691923, 253.07602567804375, 252.90375627942848, 255.8893811408232, 256.6076032965574, 256.6051837229738, NaN, NaN, 120.096037201686, 116.4474912377291, 116.02223058224439, 130.94988585898292, 176.9578761036976, 186.23833196049287, 181.4402729371609, 184.78243216455786, 196.14161111595828, 209.1555621209043, 228.59208218569304, 245.6802277537727, 253.70715658480205, 255.80705374230288, 256.1983100617013, NaN, NaN, 115.80508502197358, 113.80174646156247, 113.44228260402096, 113.40546721637564, 114.69048540078742, 131.1625345273828, 171.39634144760467, 184.55445283743427, 183.6249799821622, 199.84647885581018, 227.0280373231932, 246.05373189644084, 254.7426679104534, NaN, NaN, 113.69616816240658, 112.49678262521093, 113.05654212472005, 114.77593896730698, 114.7314296145973, 116.74136818440381, 120.80296136953122, 141.87758127411925, 176.56151561514264, 201.93849834026776, 231.4125556174941, 248.49652528932077, 256.50770331568225, 258.8498496675888, NaN, NaN, 111.79246441350757, 110.77642628386884, 111.07878315296543, 110.71865919116637, 111.6744308494111, 113.61197605284481, 114.8890687977376, 156.1081461170743, 179.39260082858434, 213.45331483049034, 238.36580909876713, 253.082278158484, 259.5026348305295, 260.47049033965857, NaN, NaN, 111.42377552473476, 110.23123700130161, 109.61795441386234, 109.29230646905702, 109.55663180314177, 117.45443498434808, 142.69920998363423, 178.17892939175027, 181.72617430292456, 179.4714832398747, 198.18737600893547, 227.97023436999862, 247.16182466747856, 259.5789751226675, NaN, NaN, 111.1362225487878, 110.30591512617228, 109.46989791556896, 109.0278406602257, 109.39716772874024, 126.33641734016177, 173.70789819997825, 188.93204766910168, 204.37538750296028, 212.01955038501183, 219.65976670054587, 229.73221686072495, 238.20560065481862, 252.7704099607414, 261.8978405054117, 263.09419771032174, NaN, NaN, 111.21906132143243, 109.73005950603067, 109.70250070887374, 109.37045176261711, 109.03602007114002, 109.28436124145536, 113.94159459471314, 150.87936264923718, 178.22114893986574, 201.03342255916, 221.9318294612232, 232.484144717815, 242.20748074877343, 253.37826661102088, 259.7382059039332, 261.20707905913724, NaN, NaN, 110.52759924719679, 109.77028838501703, 109.74275378150237, 109.70190598125271, 109.66000383430125, 109.98834764033228, 110.30782341146241, 117.61428248668096, 159.79882582826812, 180.49183695276915, 198.82229497767813, 228.0092872208664, 239.3847244499487, 244.90385950981764, 256.17082192131755, 259.4718534823933, NaN, NaN, 110.91418233374351, 110.56419533218241, 110.53371325313988, 110.4897515254368, 110.44941028192255, 110.0782654000649, 110.0385663150161, 109.69791007087086, 146.71437239330578, 177.87479583650938, 198.08758748017027, 220.97108991597784, 229.55150532543107, 237.50317217048902, 250.21748582326313, 258.5691971217811, 259.2081218534497, NaN, NaN, 110.72621533534829, 110.19125728998493, 110.16563483271287, 110.38672818322578, 109.59935623893695, 112.96904290958248, 143.53664754935448, 173.93114458005783, 177.40207866985253, 193.94943918190958, 209.41713001201825, 223.3594185124222, 233.70353840814423, 247.4155745104324, 256.1810358551155, 258.7377985765813, 259.2315376783792, NaN, NaN, 112.20294720198982, 112.18821940716778, 113.1533817336558, 113.44011607584837, 113.39908939876126, 113.02816040854935, 111.69451219283906, 109.38496211752222, 133.85587668386043, 171.92804194991365, 183.66885483584412, 195.5930311523504, 208.53114692639798, 224.51362561073714, 242.50075517822066, 255.70380221540418, NaN, NaN, 113.8294028397139, 113.5155922118242, 113.4854114406263, 113.44686339780279, 113.40800744085334, 113.66762393783196, 115.69887493516248, 117.1233824712957, 115.65906175279753, 124.45893061140306, 160.11902402157122, 194.46208945583743, 214.22331886831554, 234.08654321741844, 248.553468176115, 253.2541725900725, 254.42040806801037, 254.7024425653746, NaN, NaN, 113.49928324824477, 113.25649739350187, 113.22806273579451, 113.18870305483735, 113.14855411038747, 113.33317604507738, 113.97080880618499, 120.55160384444802, 138.35742217236844, 155.05030651519883, 160.0698019072646, 171.1392774856956, 186.579719587287, 203.9517550112238, 230.88706459327793, 250.22680860245512, 254.63178473094823, 255.27870423989125, NaN, NaN, 112.35314982584504, 111.81948702176201, 111.78957854785834, 112.26285657196983, 112.2164142909035, 113.2011143114851, 114.70476865865238, 124.43293566286928, 151.42646215566472, 170.71390635223568, 181.31545989585115, 187.81468164281833, 193.56718258758417, 206.27180022169932, 234.91782941289685, 251.25070804493797, NaN, NaN, 96.45873779167147, 99.79206565860231, 103.5312669343217, 106.1583793128764, 107.45676082807645, 108.5375396816129, 112.69597785458686, 124.79698374485922, 145.53093575174447, 168.9416906135335, 185.14035536917305, 192.01255653202827, 200.91396476817562, 209.35712086337594, 228.32125878146695, 246.29280346902098, 254.30173793144928, 255.57999669842798, 256.0038864946932, NaN, NaN, 99.4716650505386, 101.69730714568409, 104.55142110825278, 106.30049195094607, 111.80329938193914, 115.74480201227794, 128.28869244890117, 151.68002887583154, 178.71546075335982, 190.24863397589556, 200.088597736919, 209.40701403460167, 219.18360475991926, 225.5723782222384, 232.585712057542, 244.3170536251796, 257.84734892542815, 261.3722700131545, 262.0368762965567, NaN, NaN, 95.65827598816084, 97.69667235971284, 100.64898501497888, 103.7615105211178, 106.52502167575604, 107.41759714847564, 110.14969578619825, 117.46028143085506, 126.04661954719313, 132.82091468622323, 149.14476537419677, 156.81449534003178, 166.56379210429975, 184.40554511450654, 205.241714344571, 218.45929625577057, 238.95357132617903, 251.51931199245507, 259.6111792406753, 261.4213883462409, NaN, NaN, 92.10576172635245, 91.87749624488332, 92.52482922454, 94.52560926101279, 99.88188245117135, 103.42264516144552, 105.63026669588294, 110.91398183824732, 119.263558128996, 116.1632495353438, 120.13032286022863, 138.80423700465965, 163.03156450957914, 180.7254844025044, 196.3521350961562, 211.10721537952273, 233.55235170946872, 250.86632977470762, 260.69589058614275, 262.45896715009013, 262.63842615011, NaN, NaN, 96.72466105960812, 98.73510073566436, 99.82461963571677, 102.07213890236221, 104.47571049971306, 106.41913452122577, 106.8230405675792, 107.9198327100272, 109.24652189554655, 114.5632908261265, 122.70299798908384, 148.90585785058636, 176.30619868394766, 195.8764986990574, 210.22498229789957, 228.33470617211265, 246.01629975771877, 258.04290962399216, 262.41871256618197, NaN, NaN, 94.18243723653679, 95.47538406224028, 97.79797903996635, 100.63103712176448, 103.2198901980411, 105.51572201687523, 107.02887805261828, 109.34317021907162, 110.89600132442762, 113.73584696556999, 118.62252093834108, 121.96610295938585, 123.75963507184298, 136.93803326026247, 168.7271694260183, 194.68988375753364, 205.36191077936638, 215.28782698502908, 226.79102602686388, 245.8786700790386, 261.49432815819847, 265.3792625272224, 266.03719849217254, 266.22475126667536, NaN, NaN, 95.75547428201145, 97.04207117433009, 99.43542041878788, 103.12404510237813, 104.39009066149562, 106.58927628796194, 117.44677253059501, 117.06449421409161, 118.7003295990275, 126.18575295353882, 124.36170282088206, 122.20219238443168, 130.6766553738942, 146.16738136412647, 168.83988614080425, 188.91597691298415, 198.82577153266706, 209.88297295260426, 222.15934624252313, 240.15833195393998, 258.06441860801357, 265.22488369934433, 265.72132134057637, NaN, NaN, 96.87675099414527, 98.1632489325552, 99.80554012231761, 101.6455181407539, 104.95869313022364, 108.60378136404717, 110.23589096850372, 112.24308279441458, 115.36600980982762, 112.82350484892842, 111.33055287335132, 109.68304681084096, 116.48924735224657, 124.7948822590854, 141.68136832263122, 161.1836375281082, 184.2323094042495, 204.12433349537758, 221.81187501023894, 240.11382010007438, 255.78929022869949, 265.32261023854926, 267.1899121518594, 267.8522271328082, NaN, NaN, 95.97561437750802, 96.40524909327817, 99.06087065126692, 100.80607993408965, 102.1209308786783, 104.7468141881943, 106.93220524380993, 109.5627711559905, 110.9021282899608, 113.10768910187078, 115.32704742966978, 114.87734827043343, 111.37183748085636, 111.84012502049524, 115.35548706687653, 136.54771109749475, 191.10069907722553, 213.80976551477562, 223.26187929485513, 236.0198948456299, 250.91195317959662, 264.182241347164, 266.68448089650263, 266.75317712029084, NaN, NaN, 86.50986501173017, 86.87708240197462, 92.41970794231531, 97.1905433735964, 100.13682665579806, 101.9495349186032, 103.7728458337808, 107.80401124376597, 109.99412108363363, 110.7269757744453, 113.66123148593158, 116.21251016071786, 114.77191295408578, 112.29193176675977, 117.43808425509242, 143.2099849676203, 188.62836193503182, 208.9806971181685, 220.26694995414096, 230.03376344492858, 241.8548463518896, 256.5424764561295, 263.4706202116904, 265.7084642922574, 265.3953523523028, 266.16718199496506, NaN, NaN, 81.9019681416162, 81.91209427127659, 88.55710833663187, 92.59310890365239, 96.64872743495015, 100.32741920228597, 102.88140417205716, 105.06814896987512, 109.86778777397038, 113.9863592158062, 115.46248964107315, 112.15493419971233, 111.7991186071247, 119.13959558410298, 123.54569911931677, 130.53183927574742, 151.89537280739168, 194.79884291025314, 214.48082268170774, 225.76094153645778, 237.2928915329905, 250.178733677631, 262.24988262857886, 265.99378581066924, 261.7939620858285, 257.37129779946673, NaN, NaN, 86.15985393023983, 91.47211310860233, 94.11760010791441, 97.65554224843521, 101.4811265238007, 104.40950998474285, 109.70452918195366, 112.92406682182448, 113.19915639842664, 112.95618687839584, 114.12732393535052, 115.90243545549355, 115.32605350151384, 121.2087193131981, 146.2894606884232, 182.34730716841503, 204.2770818416197, 224.40064441028792, 235.83873876849813, 245.08418812316808, 256.6810030132405, 261.32540586310364, 263.0802046519512, 260.46027560223445, 254.34687793496173, NaN, NaN, 85.2266057977091, 90.84914412359656, 92.89999401286721, 94.95142685218816, 97.30271067730104, 100.23850014990057, 103.17134483095127, 106.09564101894988, 109.59958304822017, 112.81702530529749, 114.84803318558083, 113.115983155316, 114.34206433899801, 115.86516827184506, 119.97420623744901, 134.72063988183555, 168.9715363520088, 199.172926911399, 215.87535303198464, 226.37289052377923, 235.6923266823267, 248.906422953376, 255.53165203433483, 260.7718047507704, 261.23389185867086, 256.0546343139023, 254.20271945138018, NaN, NaN, 81.9462273632354, 82.27082999653315, 83.57690676983233, 85.54518661698411, 88.8373440307978, 94.11978672505218, 96.78828892352456, 97.7740136724797, 99.74768605159227, 102.04395608138138, 103.00651389788278, 107.3208309492485, 111.60274162546123, 113.2407515470191, 112.6447244858963, 111.34489340106096, 113.0420558704895, 131.60455832853205, 162.53173882011257, 200.17080516585852, 219.18744647939477, 233.61866527486538, 241.9678702908866, 249.0367462451561, 254.7095174213877, 259.7290507614347, 260.6737739902069, 259.43416539513294, 255.43354344996015, NaN, NaN, 60.58624286432823, 60.14160550258079, 62.3472715866527, 64.68558412962165, 67.16352944240353, 70.6751228698757, 74.48332992579995, 77.25355933998573, 79.1395246862936, 85.29263662131416, 99.69922142586182, 108.22213976219463, 109.41492105709655, 112.06666864152952, 111.48774318780362, 107.52006293603245, 107.63874109858817, 109.37664295596652, 111.15540482881232, 109.32278729743544, 112.15169216534971, 136.41155842974473, 173.5880966771833, 199.17123375455566, 210.55929738005133, 220.322655152643, 228.76640444246584, 240.72121855460966, 247.85665394343414, 254.18942969053558, 261.4816376142461, 260.93845484504783, 258.44986741481335, 257.81768826077695, NaN, NaN, 50.411803496361024, 49.74340252881018, 51.06664114338544, 53.2724672968504, 53.92089839385424, 54.792199679187455, 56.47769808189231, 59.34527498342529, 61.398559240074285, 63.36469719158925, 64.446204196348, 65.40098080830361, 68.1160181801223, 70.6046190238865, 73.37814434177355, 75.55506115732312, 81.34980741541393, 85.95864545778528, 94.47913718624764, 102.45985106160215, 119.4379959040532, 127.11718196952049, 131.10873614255948, 135.49526451708817, 136.5995161076378, 134.9330424192662, 132.19349387068564, 136.44202077408403, 144.3739537563837, 151.24684660635194, 163.10422712944768, 181.96925671075041, 198.30045578133058, 207.73674614813808, 221.2317409978057, 238.0794312837798, 251.4217485685309, 255.38791968284264, 260.27902687515154, 262.8599449418192, 261.0829839169048, 259.8167378329861, 259.72123717874837, 259.68299138890853, NaN, NaN, 37.79106491106618, 41.509779030721454, 42.23276075054831, 42.32849492354368, 42.31470260535552, 42.335962345688834, 42.282111240960226, 43.77834770178423, 45.31036947002365, 46.58582386657729, 48.4492454198496, 50.53255413329133, 53.56952722375467, 56.47183196183805, 58.66390718833632, 61.148579088472026, 62.78775986112792, 65.35456204010727, 69.48942824821266, 71.67471883282411, 74.09440761809012, 77.06256819181168, 79.79809446030599, 82.31523256320331, 86.95011235938101, 98.50230668957292, 106.30885483654995, 115.8497648532146, 119.68217720229633, 122.75265898803399, 126.47495648636244, 133.30706842362036, 143.3459289116195, 152.70425603872135, 161.10682065599366, 163.8805427424063, 167.4566532401184, 170.85591311532423, 175.76115773799742, 181.23202945727738, 189.0556665861956, 196.97585331702334, 210.53956978961978, 229.23110284470314, 244.23046612407154, 250.95581740554348, 254.15088190936697, 261.5910651428647, 266.9053641163907, 263.5433471644329, 258.88009097118197, 258.3690383916466, 258.62995537053087, NaN, NaN, 22.98928504191666, 23.02666382659477, 23.72258328000363, 24.49029362698323, 24.924833189067474, 26.099877213489922, 27.126804937615052, 27.968331371620067, 29.954084750895586, 32.1570227709789, 34.4307917099012, 36.22241880402378, 37.24058261238052, 38.076542233960424, 39.46545015899328, 40.448185595398975, 41.986769932333765, 43.96766180772672, 45.28257693280282, 46.52277009161366, 48.31654446464977, 50.51379110983057, 52.637121368501546, 54.104176294685075, 55.4916397660924, 58.27442906385698, 63.40390397199616, 69.48786981986714, 74.4661043039604, 82.60439517507677, 90.14953328814755, 96.01584601150088, 97.25559565923359, 100.4735301570803, 103.47648207027741, 106.83611945976168, 109.24133274544694, 111.86558019436484, 117.5731461017002, 126.08306971261848, 132.9549417587016, 139.86075520834186, 140.8840620349316, 140.42761234630734, 140.55856693705047, 143.7958575723362, 147.21099063399956, 151.3325014450337, 156.69494717918457, 163.6891587696977, 170.6664215118262, 178.23838079119395, 182.50687076353503, 189.1115864397851, 195.40040721755017, 211.942944606653, 225.45070276922726, 232.71473352323278, 238.88762635059715, 243.74719308346172, 248.41036264135644, 251.9729580081735, 254.34316277509942, 260.96688434652356, 263.6151306690939, 258.51126626570465, 257.8725771131952, 258.1204901948345, NaN, NaN, 19.994228084467196, 21.17304138555189, 21.61036600378389, 21.749102938546127, 22.482098463247276, 23.36395746984147, 23.432969645180222, 23.35556204226979, 24.010523579339832, 24.886025323724997, 26.132018931145254, 27.59675253394622, 28.61873650920407, 30.00799111146262, 31.250615680444746, 32.56566468234876, 34.98390319027787, 37.987859306438395, 44.738005041865115, 48.91478358786037, 55.80601214950849, 60.56853426462462, 64.08352198155174, 65.83662191618899, 68.02970983347106, 70.00560901420799, 73.60396289861619, 77.64806178920743, 83.30406606180013, 88.79625852002461, 90.83602386062354, 95.8132948137039, 100.42269223214163, 104.15469443839419, 109.12338264099563, 111.6761451764084, 113.57523393482772, 120.45340201496094, 125.8511936477539, 128.56107380915424, 134.87341730749995, 138.5131760843304, 139.18305781600452, 140.82888186013665, 144.93038431875814, 148.4850269561166, 152.63724563763103, 160.77146318661408, 167.7564276096491, 173.2214269642865, 178.9890387153588, 188.07090442863716, 201.68596840734895, 207.21527149864903, 214.63765786200955, 222.24034824503164, 227.6616386685026, 239.91571242260164, 246.51110995935218, 252.52542324008667, 255.7900395615492, 258.10185127334057, 263.7283384506408, 267.2223537472576, 266.07289199024734, 262.31116494620227, 260.03539365678034, 259.53943753568694, NaN, NaN, 18.077461735962938, 17.77907207535235, 17.92255615556532, 18.360334291931537, 19.091606273460666, 20.11657753237387, 21.36387624248071, 23.127625224103237, 23.85973879725498, 24.51733895066034, 25.320936732866915, 26.494053679810502, 27.442720069281783, 28.833387535008285, 31.10667821837768, 34.18821408560403, 36.97209208872346, 39.608908111127796, 45.39743491470969, 53.31803591745875, 57.782873502005835, 61.00299597928251, 65.17924739902884, 69.86695667052838, 78.07724345805326, 83.20362188420611, 86.86925884728993, 89.58630424468015, 91.27158665602202, 97.71162949677499, 99.3063584563537, 101.93601401672314, 104.50775863198852, 105.82558535398792, 106.61399060932973, 108.73095179916776, 112.23584764229138, 117.07406806126248, 120.1301995947393, 124.95767141776764, 130.2544349664843, 135.3924197311226, 135.53614192661487, 135.41266491137796, 137.60519468685106, 139.40360340134487, 146.34649777130963, 154.00580924726933, 158.88079761701636, 163.60411517203258, 170.4286378748178, 181.29963565847368, 194.64186914858874, 201.98234782268102, 203.84278701182728, 215.23707845830546, 233.17430560590543, 238.67575052375568, 242.75482446360536, 249.66126844255547, 256.5658995673007, 262.38434577932657, 264.9170362037944, 264.4098164485703, 262.27564128370796, 261.51262632656267, 261.6483274862608, NaN, NaN, 17.817770323492248, 17.70465951434721, 17.148137922562153, 17.14210597146686, 17.801209395978727, 19.013418985968517, 20.443805043758633, 21.32178862413064, 21.75857353881685, 22.85692813628646, 23.623770694054997, 24.94279591545714, 27.25593110565992, 31.107872375528185, 43.1078346686101, 48.717899863309604, 51.90626720926291, 55.53017640457608, 58.821126529052634, 62.114281661528985, 64.81954704814592, 65.98561044259328, 72.36178486156719, 79.10618807312946, 78.81289492660656, 78.29018752994077, 85.53664204356392, 91.03638118924786, 93.7452295048413, 94.89866887784211, 96.72307182977826, 99.71830235420354, 101.45456230648412, 102.77049255751744, 105.1996224815596, 111.59901124367016, 116.7955639372484, 119.13285418633438, 122.1403256835627, 120.51215691001708, 121.76933643070369, 125.41614205696041, 132.1807118790406, 134.07777679961117, 138.9395629524222, 141.0092404412656, 142.79235453643784, 146.91867235084786, 150.87456928386106, 158.22553113200422, 167.1003272695437, 179.99297138893343, 185.87953450870734, 190.74249048321332, 192.28465752690835, 200.63072257349157, 218.21593019503035, 230.94009451871173, 241.42180351519764, 250.14335880054242, 255.5720157022735, 259.6897673625012, 264.3013146398439, 266.0345209474572, 265.1187458783288, 261.89903369371643, 261.1881189059119, NaN, NaN, 20.437017828434026, 19.846637485073135, 19.109644156345972, 19.252137205116387, 19.614441797317955, 20.05221714590226, 21.152678301695097, 22.179548602543466, 22.835402626829467, 25.18312109875031, 30.104236080802, 34.290057128662404, 42.29546581224079, 47.86965430166457, 52.41771525678134, 54.61063817699241, 55.77508500762, 58.553095214303035, 62.3615633911392, 64.19681302892234, 62.61252718761605, 65.39554973258242, 68.98169219185549, 74.18220263677141, 78.06152309561526, 83.18298564387409, 87.35576050655925, 88.44216276005233, 87.55021504579457, 87.47336632960055, 92.96319237223399, 96.54640684725, 97.71074284144197, 99.68995429253486, 102.32562846357375, 106.7880093277605, 109.12440148157775, 110.51406404402586, 111.02522191947358, 114.2374291693767, 123.87591837917806, 129.60393837487254, 129.58967766393778, 130.62797185866924, 139.16607302853456, 149.89295070630033, 153.6354347467833, 159.82886183030644, 168.80128346781802, 172.19775810043868, 175.7575531351213, 179.94009061395758, 181.76466100560035, 182.7269799747142, 184.78561418974064, 193.192232524101, 203.04328411732175, 208.96003095224418, 215.20009715811327, 232.30386876405473, 243.34323657011706, 252.62274550492856, 260.0070281456115, 264.5337520986333, 266.82473570949315, 267.39006149548095, 267.2881107874684, 267.4093509315415, 267.23318551696815, NaN, NaN, 19.555687903445975, 18.52112437852218, 18.81227383668425, 19.17396533935397, 19.68415568827487, 20.56351210921524, 22.176786234018152, 25.259124137230167, 30.178582113816045, 32.155245421932435, 36.2626309574238, 42.93940279555839, 47.77800587542428, 50.929606750470775, 53.93960300375639, 53.27587516135873, 51.72661364848849, 57.36672092394819, 61.7680491555204, 65.2070078404432, 66.77371521140996, 66.91425996788126, 67.49645816345195, 69.46813576633046, 72.90672649139161, 76.7123799269132, 82.5670731597109, 88.78700457435303, 89.95755918162425, 91.9435496157175, 98.19421250603706, 100.01966705101036, 104.05234010717041, 108.14892572064632, 114.23895247414154, 119.65728382386816, 123.24787664060396, 122.36028880169347, 122.49967675656309, 124.40722282975679, 134.19604643626298, 149.45636393120256, 152.13808989673706, 156.5802391392412, 163.04323297862376, 164.20942881130557, 168.5018593638637, 174.16327721710036, 171.40659164806763, 167.5685780255098, 167.51847237377734, 172.30040646401065, 180.36395494625125, 191.11855608192377, 203.0951138299967, 215.74978207145588, 223.17695482563164, 231.57009834613405, 240.59637671608826, 246.0525415253988, 252.16540569266792, 255.32056777707052, 259.1135438043069, 262.9087755358091, 265.9816725469025, 266.8441944361209, 264.42323360833194, NaN, NaN, 19.325725620044548, 17.776645676245465, 17.625488674114223, 18.28406724585931, 20.12081298504085, 23.49739802751039, 27.612987323106758, 31.502775163450863, 34.145346225270316, 39.207750056139844, 43.16945797734447, 45.8062396452747, 45.139671263052925, 43.59669319079863, 43.66485922507632, 45.63995196092451, 47.76167370632685, 47.762274124552846, 48.41823921423621, 49.436848811772045, 49.5722294302103, 55.5095428702365, 60.71450504763685, 67.97011241131669, 75.96883468913522, 78.52587939343466, 80.05650598471111, 84.88654329345574, 87.82801058706035, 89.65368627822858, 93.53609722970859, 97.34399279239327, 100.48943355437792, 103.12378847253011, 104.86979015966922, 106.09708212832018, 108.4375398943207, 112.84319991392094, 118.62059034213821, 120.37230767199325, 126.29906602757056, 143.70507566486975, 153.80628799509216, 152.91886853427226, 153.08716805235466, 161.6150073175391, 159.8584371793491, 161.52074161881674, 167.41980580420721, 169.68407825524196, 162.24542699804792, 157.02146112140917, 160.7632460082802, 169.83229166814854, 180.77575438354503, 192.40327938671734, 203.7832783035687, 214.76459642283538, 220.72124574072075, 227.60427888755433, 233.27176072524983, 241.9047420823481, 247.23630172984008, 253.2936210504864, 256.7596493226777, 262.4546868477158, 265.17203579725617, 264.2899189384848, 262.25050006739895, 261.89736854861707, NaN, NaN, 17.408373810768133, 16.19020261744697, 19.05793322484715, 28.32548702346512, 31.744621605694913, 34.939065199338835, 37.36045476328564, 39.008241465582365, 38.234343596043274, 38.12150853448484, 39.438074906317034, 40.08762662886389, 40.96376122027687, 42.281532183544954, 43.92756182709091, 45.46058115220041, 45.23411105636367, 46.76563687730105, 53.3626326162219, 57.97449308435608, 60.01287241888959, 65.58041446630092, 73.05708009182534, 77.5955230770241, 80.5313372214534, 82.86889198179533, 85.21723152873265, 89.91015589620172, 92.67303828270427, 94.8549200203046, 98.65635256298752, 101.12756812564228, 101.98533750713813, 101.67774301914937, 103.42293525749952, 105.89756257698744, 109.41478080093272, 113.50212406127824, 126.37402728909295, 144.686558704593, 151.16164062084354, 151.77699353296282, 149.16987563777948, 154.31009413967377, 162.81905279401494, 166.55890904538435, 161.17834903260174, 153.17182555134488, 151.1760651840891, 164.22063106323412, 177.5073185823194, 189.16118624321228, 205.44024064985737, 216.26415657238311, 223.70337670220118, 229.55653603689234, 240.05779576920418, 244.80956045418, 249.46807187041577, 257.2919426657304, 262.5116104704565, 263.3160074508061, 258.5042694608677, 254.46810147153897, 254.36524648841126, NaN, NaN, 26.863168797786493, 26.270246125985537, 28.10715815114358, 28.253456445416607, 27.22185612895259, 25.305537959306545, 23.754249170537168, 26.173570758869865, 28.960239415148465, 30.421553395622745, 32.25290221636219, 34.67708899646007, 35.26047275922804, 36.14065080896041, 37.092466303568244, 38.91884868258619, 39.13539903646452, 39.64234293315277, 42.93963324285317, 47.627198877550086, 49.89026110781744, 53.10691569682067, 58.81795313255283, 65.56231287234628, 68.64465518582752, 73.03803622544797, 78.60796577063641, 83.59627088476581, 86.2252269996402, 88.71901363786714, 87.68503635730131, 88.11851104938121, 93.66946886665461, 96.73214190860588, 100.2427823951097, 104.77516993265512, 113.12926650352377, 128.66440996958704, 146.68109611911925, 152.68319246513298, 153.94738238310822, 155.98842850485633, 156.4346151799793, 152.7898203989202, 154.70703359454384, 164.0753509543747, 160.75417537141666, 158.4276212811271, 151.15581731132346, 156.96273680008255, 171.03771687173654, 176.42300979928896, 185.39288354038277, 192.96605806017564, 199.97334622015794, 209.9494980556333, 225.58269989819527, 235.25825362107645, 243.8864704303836, 254.43669890447416, 261.30882818518495, 262.85771444279305, 258.29637156574796, 256.26090238115165, 255.02555532898197, 254.19560366247575, 254.01448328921612, NaN, NaN, 21.936790747393363, 19.135086029853397, 17.952402384231007, 18.168631080524154, 20.446719719078512, 22.355505467709566, 24.264302657964837, 27.127264248697415, 28.44490440008149, 30.056120910001514, 30.274365462708186, 30.709648437663272, 33.05536910473349, 34.29863008157597, 35.03042313313698, 36.27637861081139, 38.545000999370224, 44.04514458754362, 49.62209758336312, 54.09131559357445, 61.74798969736433, 64.93197740770391, 67.67793594236952, 69.76816944353388, 74.83213787787783, 74.3931383134481, 76.15313710929064, 82.855950968833, 89.67272607410105, 93.18427689849213, 93.93890298737237, 94.9150426726486, 97.87615258373052, 101.70761837980866, 111.69447214874525, 117.62381133389103, 127.85115430430113, 125.74584829136579, 120.24262489703493, 128.92089398983, 140.43622853958078, 148.49187664100737, 158.60808225743367, 164.48235996943117, 167.0092172214902, 168.93003208387253, 162.98069599038973, 159.44976114733817, 158.8948755380214, 159.54060917262998, 156.83630961708369, 165.91443779110966, 174.7610677233503, 186.8625077087548, 203.26085477405093, 210.95561400684272, 220.11852574598026, 226.4749092145804, 232.12415088023667, 239.37813943787145, 245.97776281369082, 253.59821606730478, 258.93462337207615, 261.05881747136283, 263.74550995519775, 261.80885091375853, 256.6520686684591, 253.97212764405498, 254.22172607285754, 254.5586948953846, NaN, NaN, 20.911942344889486, 20.467240865045994, 20.906058848932027, 22.51970602572533, 26.560186141681612, 28.769429371686474, 29.352472302158255, 30.38011845600362, 30.740627816702034, 31.031072886448207, 31.90738758380187, 33.52170565775604, 36.38637491468262, 41.37800843141331, 47.981509249029536, 52.16119208539931, 55.31251324733544, 57.50828585717013, 61.01917173039934, 63.87407758992004, 65.22068433136026, 65.07223160744573, 69.76688918803673, 73.35887716483357, 78.70519156358448, 84.56795272978448, 85.64872933632115, 87.8359684310977, 87.24424599650064, 87.22816293439746, 90.14187389385778, 93.64069692305749, 94.9556849650508, 98.39356840271752, 97.0645746285563, 94.42274313217719, 101.52066860633438, 107.73860001246929, 111.25414227470368, 114.84635065756572, 135.94649358368343, 153.2348818714388, 157.92229776431304, 160.10454736999915, 165.38078316677044, 168.45739259552735, 167.31252881532566, 163.36010546911896, 154.20493599002347, 158.21878773535275, 158.98885135720275, 159.3563486348416, 165.9354897632724, 167.73597561049414, 173.8659941620413, 180.10177712758104, 185.7400978684904, 200.38464909049918, 211.8960059277202, 217.06391336454018, 227.75420879100935, 236.55518014127412, 247.64005787412168, 252.49165282201398, 257.47814454480266, 261.6902856814332, 263.9256265722284, 267.2247931536451, 264.81717076088654, 257.80363214414405, 256.088017385557, NaN, NaN, 18.44200376667598, 19.911834836081873, 21.159995241343537, 21.743864858669603, 23.72435897443323, 23.644647674104313, 24.81500783830369, 26.86907805199335, 28.703388489700085, 29.436323545699732, 29.79693949338117, 29.937389658622067, 31.39951575328877, 35.507876491261804, 41.1577797717901, 46.95165243669177, 53.70294358200689, 58.10102356804552, 59.266391718502454, 58.95764468548973, 59.9028010858722, 61.989176480798946, 65.72605368488458, 70.00861133707198, 71.9874269143174, 72.8659463083905, 77.03881478853364, 81.32494677339679, 86.59072805779054, 88.23081948332974, 89.31725522597787, 89.75466164004884, 92.061499731171, 97.54903484169141, 101.71257695605458, 109.29559808721645, 113.7953569469164, 122.13312773217297, 132.2568232902426, 144.0059386244071, 157.51373936558485, 163.9492853589992, 164.8186601916345, 163.08631711486711, 158.0024323657651, 157.78204431113693, 159.71140720381695, 160.02891533947349, 160.3924166048793, 162.6525039435018, 166.411844051944, 171.6694162754696, 178.81141770543343, 185.21186177889382, 193.67048431539874, 201.4379619274198, 210.87204157066105, 227.00756378939082, 239.83054291162077, 244.97530442521648, 249.24848027341483, 256.6085739163776, 262.37466636595616, 266.2942134489902, 268.1325936710377, 268.9640315410721, 269.1932674003688, 269.44325814098517, NaN, NaN, 19.76022028633627, 19.168014931178945, 19.090657385429783, 19.23190689055158, 20.036739904116843, 20.987474540365458, 22.159766438100636, 24.652565694803062, 26.265118853931394, 27.071084444583523, 28.24368905242679, 33.52655628550458, 41.086344017329274, 42.55432517668324, 44.60522453203887, 46.95162219975613, 49.15060276387215, 52.007099880392865, 54.49646150197034, 55.51523134609172, 59.32280716008051, 60.92287416048959, 61.64755970672468, 64.13405660816524, 68.83244429718722, 67.07947527514908, 75.80158743069065, 84.74046301547462, 88.32781390533896, 85.02577138681258, 85.44860951345697, 87.78577769397535, 91.22899429678405, 96.8610649781761, 99.0479582170035, 105.04355553406945, 109.07242416541058, 114.55957202904078, 118.36061834866739, 124.20695009175252, 145.32857919903086, 158.0649086604552, 163.44701214597, 162.92439806529757, 159.085020692257, 155.8105466981337, 153.53066272052482, 160.67672234977414, 160.76526232287495, 157.18568273190533, 158.21754504689102, 166.00905242877658, 173.9979601057468, 184.1865085436596, 194.68896136503156, 203.6454488673082, 215.64000982785262, 229.28813544520054, 237.757756678942, 244.0180980908798, 250.57956740728025, 259.2704163121833, 264.46026334276087, 266.1869467743704, 266.1361342318611, 265.9547736564398, 265.8352167988587, 266.0055082467381, NaN, NaN, 19.725515140602273, 19.022758364297818, 19.791961022370444, 21.55521969250761, 24.424425758982196, 27.656523434955915, 32.09934956217541, 36.395157190113196, 37.30782988355122, 37.45167964159753, 39.54237527378658, 42.445049422325525, 43.247368415354515, 44.63994252783065, 44.77765170706371, 47.599910535594425, 51.891499913758516, 54.74697632864204, 56.396071345018214, 60.23660871717337, 63.7167133969825, 64.6672871338591, 63.335019397241666, 62.01049627265981, 63.09983260243249, 67.92752836018481, 74.0073071855704, 80.74562835811163, 82.93944152301701, 86.23471356054601, 86.30142759192663, 84.46898368934329, 86.14644224503861, 93.46469669688986, 97.63480768630896, 99.08711147392627, 104.49482101214694, 108.08055441870238, 110.78666000561516, 116.71435586876176, 128.1028490475765, 145.10097229321084, 156.5205364815829, 161.64681925772766, 155.07096291351178, 146.9962671650879, 152.706652065068, 156.4698956375187, 159.176603597614, 158.03084693257887, 156.18387096016806, 160.19490999290667, 166.11770327628506, 172.56268349129363, 181.4240650752831, 193.03780347260948, 200.71289981168232, 211.69506423417423, 226.19205768871237, 235.0437389632932, 243.49439880195672, 249.87254497010682, 254.82438883647984, 259.89689668761184, 265.85319538013204, 268.3551496878065, 262.5303455749569, 257.05795340893, 256.0605608157305, 256.025658410394, 256.0750656853912, NaN, NaN, 22.751674942190323, 22.52995924272087, 24.146982437332884, 27.820009485373497, 33.48494597764121, 35.02703923243889, 35.68077461378684, 39.20238989230231, 40.07398741145922, 40.43706857580446, 42.33827477551183, 41.88797355793053, 42.68869747294307, 44.29991369417539, 48.189235424549615, 52.810194226815156, 55.88601295028086, 57.48924934827779, 55.937094387971314, 54.75355155690135, 57.7155206008775, 61.23129539792375, 62.43732972704733, 68.16013592239426, 74.86629196896006, 77.61133324381467, 79.80468964176414, 81.6602685779282, 82.75427023347041, 81.10387066138311, 81.31435654720504, 80.31546541711322, 87.78191328210386, 93.60122909218339, 98.09174418159597, 99.29537463369792, 107.0931641256152, 108.9584055549634, 115.87339040627565, 126.08359553119334, 131.16866631482193, 142.8820890992003, 151.97537817423452, 159.5983112789075, 163.11071151236303, 161.3280152064995, 146.6965311592338, 151.2825484396777, 158.05578446403732, 162.69342737165945, 161.13336657143634, 159.35153154790734, 161.16177896792547, 166.51238360156788, 171.96157205243702, 188.73001844416976, 202.63560447152085, 212.61362854415685, 220.6712161037255, 226.36770947012275, 232.88070514214226, 237.90249283817613, 244.32975617624027, 249.3917829457555, 255.50825155683083, 260.79109822963073, 263.2421101537409, 266.0436490007714, 267.9843247842508, 266.2526141596187, 258.2120326853015, 253.7428618618724, NaN, NaN, 20.645803338617792, 21.084931615659947, 23.47600644538799, 25.971571707080106, 29.09380416259793, 32.36152995356286, 36.43852158157103, 37.348912826751466, 37.52328925648296, 38.251767211022766, 40.415412054346966, 43.46240185678998, 45.5506431815662, 46.68149733963309, 47.297474254268096, 49.71043464229692, 51.72317606190617, 54.39722596836566, 55.233409246917766, 58.15741929628989, 61.48838799667513, 64.42061485683129, 67.49663950299932, 72.33037079707111, 76.58484801152841, 78.04339080806194, 79.21374597593898, 78.3311188308464, 77.29529784393651, 82.71123103157358, 97.07037313328757, 103.3739925695043, 106.29576612130352, 108.03974261259329, 113.60515727560302, 128.69660451816264, 132.06189421073432, 134.39897096098596, 141.4285093195704, 151.09425456873106, 155.66089912473123, 160.9442568641849, 155.91023416481903, 145.35775219110315, 147.84992152746113, 150.37718538485075, 145.60971960027638, 159.21401866646312, 160.68591609608742, 161.16412634231344, 163.72515322821496, 163.9748219138592, 166.15351493107218, 171.7224573052969, 177.5588832301173, 183.26950068276835, 191.7121132718259, 198.61251846917443, 206.3726135815778, 210.7639512784606, 215.20476696213206, 224.91670275709677, 234.24841735431608, 240.98052493006418, 246.80010045243, 252.70440539149982, 254.6971516974208, 257.30488215268133, 262.13003879515276, 264.6538524882761, 266.80015017440036, 267.3045268344837, 268.8341540913818, 262.24346438262256, 260.79329174306804, NaN, NaN, 21.30837478088452, 21.010753957036453, 22.553244918236373, 23.504586591894476, 26.66416812677908, 30.853868811536852, 34.23344489609096, 36.14355114880908, 38.04630928768127, 37.3793731940628, 37.220116141608884, 38.45915277687526, 42.34919089302731, 48.07489362935766, 52.84338404713766, 55.111815188300234, 55.46880639990142, 54.57965650358648, 55.822051173339936, 56.68834004146912, 58.07239946296888, 61.370730385391866, 64.22623138764226, 67.29853842169638, 72.57549247961754, 75.97775511290845, 78.05920294967554, 79.3729057879062, 77.93415875243721, 77.49112542112779, 81.77074192404672, 93.4170915034611, 102.09452523633479, 102.74468797659502, 109.68101168368874, 115.93564081011868, 124.16748158037315, 125.81239503025105, 127.65543478959343, 134.3589704574862, 147.85143531332417, 149.1703129442471, 138.91467302782016, 140.3706356659279, 147.5294021575358, 152.94694637202568, 147.38481821685053, 141.68231365323695, 142.71282658816264, 157.44205814903856, 161.9738268574944, 161.54760461525802, 161.76802529883167, 166.39455722690553, 175.34721699141937, 187.66119420947766, 197.39677023099625, 206.2226267461019, 217.1741839302331, 226.91543591651623, 233.43039874994938, 242.74081349276364, 249.29043172493542, 254.42562248226133, 265.5514230657701, 271.09894639361715, 271.786213894596, 266.43426314750906, 262.877439345136, NaN, NaN, 22.560486634760288, 22.85101962727863, 24.688309074359104, 26.228979678919032, 30.124772849850743, 31.66239742992006, 32.539148517269666, 32.38814901747673, 32.59970505204361, 35.8988277184879, 39.41341989323497, 41.01971925421735, 46.31033664084934, 50.562699888788565, 51.87690691399318, 50.036116687810235, 50.172941104525904, 53.32091628570008, 57.79308464174615, 61.16094960272587, 64.52610072467053, 66.82779109338529, 68.137107336525, 71.32045768028121, 75.71528527750657, 76.70324262604385, 77.69083320647601, 87.68856334143877, 92.40985521505948, 91.73984766630683, 96.66941064358141, 104.36418596345864, 112.72644187166641, 117.8897504871977, 123.80980678448906, 128.7418610576686, 137.430566091301, 136.21781223511957, 132.69102504623234, 137.08198767844286, 138.97127944597736, 136.32743924825428, 137.92854728526862, 142.3058249923994, 143.3400535619827, 145.25624341663803, 159.05243534837751, 163.82120976503774, 161.44572814692845, 157.95041461261806, 157.25036914285698, 162.01028041933145, 171.70660315329224, 183.93873135463826, 196.68487721425612, 207.62475202461516, 221.86941698955766, 230.84229356834695, 239.56812895795994, 244.73556721958587, 249.16680819158813, 252.81608256205539, 257.0225251516278, 262.3536545095845, 263.66471226604597, 263.90395812714735, 265.42872082785055, 266.13631462334763, NaN, NaN, 27.670958662080878, 28.182198316525348, 28.471959751713165, 28.836490285015056, 31.035803119728406, 33.97217396745406, 36.099672096447684, 37.04327028220027, 38.28397938879627, 41.731995043349244, 43.55834080767911, 47.00581397755577, 45.016753835976466, 43.46865509270692, 46.030767593456154, 49.39952876293645, 52.18418282147434, 52.47467585994193, 55.108263044223136, 60.170386511166164, 62.69770836718659, 65.04202574189385, 71.06103658922413, 74.72385216761073, 76.26652345905516, 82.72175663782713, 87.69680461337606, 93.33633989980999, 97.21292156712633, 103.14266348409738, 107.54164644932915, 115.74862604026889, 120.13453365693928, 124.22963873303271, 127.31131586747357, 128.25610315499375, 126.4834272571066, 127.20509954362227, 128.43393189977252, 129.08538603441403, 133.04711069555267, 147.41241766778012, 156.48164889405575, 162.92119702353497, 162.3323036355875, 146.9896724547559, 152.5687397662772, 160.9634974858161, 161.7534142774872, 159.2842107667765, 161.08503925150578, 167.529481203671, 178.72968397603293, 187.8718677605342, 197.45352594779663, 205.79327660722308, 210.41767348915226, 217.783577320316, 226.3259190403357, 237.58956749729583, 244.43072100503466, 251.08079515128324, 255.7937068886979, 262.84046327993246, 268.56110258971836, 270.03018337413977, 270.3182007092356, 268.8563041272156, 263.0425971896957, 260.7689073791145, NaN, NaN, 30.369229902328037, 30.142913250506474, 31.391544605211664, 32.19379109383738, 33.65775231777573, 36.301362064875605, 37.39658604492023, 37.532048877837816, 37.96699679096726, 38.769651063599795, 40.01096145248848, 41.99102946299535, 44.26500093586458, 46.826609464354206, 50.71408829454575, 51.073535379780445, 53.70476677895066, 58.83601727181591, 60.88486329206799, 61.98095755777767, 63.47978542662582, 70.62301798520967, 74.24515343846561, 76.1069033834821, 78.8536724095772, 82.81542814614764, 91.3797903414436, 102.03384836852852, 106.20968011229552, 106.09519458998643, 106.29597613411086, 113.54559334458243, 118.38471555091132, 124.63629122474298, 131.65358234552832, 132.51532510090078, 129.21163649729414, 128.00772942175092, 123.61342195286107, 124.165405426005, 130.4925164048311, 138.69634132624557, 138.69255769821171, 143.82748940591682, 159.06689684182257, 161.7300034710655, 163.94535782913505, 162.98513056065823, 160.29103669528666, 162.2026346687503, 167.27074747212495, 171.8930685451687, 178.02458457162945, 182.37833742437115, 189.84094954922995, 196.06452144128423, 201.60809058733673, 211.18966492678348, 225.26920525744814, 235.75251711971296, 242.94746535142264, 250.0844179702474, 257.5318326741646, 261.54038615154906, 262.67546151107325, 258.1142045720638, 255.6358202027029, 255.75025043024954, NaN, NaN, 28.4111291917869, 28.481881998263454, 29.50778342091554, 31.638139232459196, 32.95735212208016, 35.0132518910864, 36.623044381008484, 38.74927769050149, 41.53569700589202, 45.130913083366686, 48.28758327023546, 45.861279925897726, 44.601990948811995, 46.13210927297886, 52.07265241518702, 54.49102241670306, 56.32307687194859, 59.18645770502272, 61.74541785830362, 62.984128092275114, 65.725539613492, 69.09195417517212, 71.72652384353388, 73.25612065067824, 73.3992288228399, 76.69033151343042, 81.15275710705069, 85.1668335183667, 88.89468610537195, 97.16748689990679, 103.31386568257979, 106.83173238011841, 112.25494347011222, 116.84542926131343, 118.35959961240668, 123.41097114048885, 130.37066100213886, 129.11434770800028, 128.1647832188038, 126.85393139081434, 125.67314579036025, 129.46824344872977, 138.86868048357596, 155.14175356055728, 145.33868061614731, 141.96278908049308, 160.02532273088457, 163.70509376410064, 159.27200369407427, 154.3601885241602, 158.09413304400658, 164.01342781684215, 171.56872234588857, 180.1968511321799, 191.11838126009204, 197.69035219245632, 204.0999293142491, 213.20020208323245, 220.48002591026577, 229.27609963072538, 237.28887514214486, 244.3957376502793, 253.60768864533972, 259.71993731524253, 262.17714005110815, 263.9664346808993, 259.5475513726796, 257.41994974411233, NaN, NaN, 26.489761104907455, 26.044716907212244, 27.108809986707794, 28.75833011078322, 30.297428700071983, 31.726356059623605, 33.55694739806276, 35.977674724041705, 37.62475707482788, 39.898755418292744, 42.53866824941966, 44.51583591474623, 42.27090833691777, 42.92393603222219, 45.62990803021451, 47.236987115412965, 50.569667156715106, 53.7603258930476, 56.50256596375623, 58.58581767325128, 59.71666581765499, 61.32158282890247, 65.56652161178812, 69.59223071965823, 70.39263076276308, 69.80127590560667, 72.35679656976156, 77.17865110538146, 80.68811472895997, 85.22349277608836, 89.97319957311679, 96.85633002813097, 102.71105133985787, 103.87886734148626, 109.29217257093116, 117.10995980522783, 120.7730846161344, 121.66994483122903, 121.38593820630744, 120.57114385290832, 123.7196396417262, 125.0502398235439, 133.08754208474298, 139.45363256718727, 141.55242139370245, 154.63271666467983, 162.2479282323077, 165.23200178267604, 160.89627021476178, 155.1216172915889, 147.65231980376493, 152.20395751406068, 160.75874653770975, 167.85266034935367, 174.6332910231063, 181.99013548844306, 188.66903115685162, 195.70683816655793, 206.7435481259569, 216.48038609600675, 225.3832472880662, 240.06140453436336, 246.9840606075849, 258.1056128986913, 267.2965978154971, 269.66478324342063, 269.2059892154883, 266.93156021649554, 264.96971572284207, 263.7563113920904, 263.8723414619197, NaN, NaN, 28.29848611143069, 27.669418661785084, 28.51085028693576, 30.308008188138896, 31.699132944070037, 32.650086775922404, 35.440505985607224, 37.64212482336552, 38.703292484689044, 37.63263278077229, 37.58528940097434, 38.38809457121213, 40.18223311004613, 42.6334776319827, 46.22408092688994, 50.18182902381767, 52.858522063072236, 54.06258012051406, 58.23827287733601, 59.84132121035987, 61.15792344847209, 64.8948414686475, 68.07944742816731, 67.19676242310501, 69.27508627501119, 73.6644193716938, 78.8245835676406, 84.31694696855897, 89.68836454075037, 94.51967679317123, 96.48385195546932, 100.21779140696582, 110.97938822877717, 116.02161260448216, 112.7170214952507, 108.96663951698704, 110.29032931099381, 122.39147690498206, 124.82086116193936, 125.7969495423067, 131.63012163874114, 132.84664452652558, 143.74571527715813, 157.1671428242705, 165.41371257135674, 158.44166892538325, 155.01672500057694, 155.2435068124341, 158.8485316656579, 168.56498896704284, 180.3262355055005, 192.83436521051243, 201.5740306276752, 211.6292122490304, 218.68986527238727, 227.9283408319399, 238.40769657033886, 244.43336402283714, 252.43578700542378, 256.0857703735901, 258.36856896075665, 261.38889562869684, 265.914349634358, 265.4065560614275, 264.9036425427536, 261.5525189783372, 259.3605686489393, NaN, NaN, 29.408365941960188, 29.773287914854453, 30.57896198724855, 31.233948948177847, 32.40358574495555, 35.04666600963796, 36.14220566460233, 36.50326559269571, 36.86516847845489, 36.712223110263544, 37.58788581325696, 38.09493934746805, 41.3228093172065, 45.28316105124849, 50.19546754539162, 53.71221889048362, 55.839865393549424, 56.34568512515645, 57.6580868908169, 59.85465395261985, 62.67000079759087, 67.14649335469353, 71.5446067470436, 73.74354639858714, 77.83972684948205, 83.33217472171054, 90.1462569813785, 92.70701844142386, 95.12856090315964, 98.56410414863393, 105.38164812331067, 112.7639914659865, 116.04469236100498, 113.18399812099705, 116.09438870719498, 114.45848934957941, 114.96414811797328, 117.23597421348289, 115.40412759115823, 118.39147331721051, 122.78334189901656, 127.74500944189278, 140.5707612781197, 159.99549661952028, 163.86644677660226, 157.68565777678742, 151.86658170907364, 152.61907530749576, 155.94228695963477, 156.40477693680475, 162.5151729056456, 172.75292414496846, 183.4321146957995, 192.156088412044, 202.38058291091292, 211.765394663616, 216.8242352042268, 218.66188601843038, 221.71601923348848, 230.5740319295998, 238.29095161252394, 252.44377894846417, 259.41973299861195, 258.7051501632273, 262.4484578139835, 268.3924529915705, 268.43139681073364, 265.5096303429311, NaN, NaN, 30.517268732101822, 29.55437196018902, 30.692100668455343, 33.445815678993895, 34.76188414967941, 35.5656518739992, 35.414320800964596, 36.107558215675894, 36.87203084206315, 37.968803576807964, 42.1145229596226, 45.929568157385056, 50.038182551257755, 51.17512831188155, 51.46224971454108, 53.73283479350496, 57.46870374134437, 61.32332736664941, 64.76986572127257, 67.91771650673334, 73.55435638434923, 78.82390682508532, 82.33146738255611, 87.93557874860203, 90.13041323117184, 90.11975838131202, 94.07126925807574, 98.13741052453801, 102.53870916344165, 107.35753530995333, 112.73607577548565, 114.81523998530494, 110.9508086570727, 108.85846116188007, 112.37755966647983, 110.28120396671495, 111.69567541032067, 119.48151229921008, 122.67324234414735, 134.88646924224176, 154.043189498846, 162.26111908306896, 165.53584330234818, 166.32046845046187, 163.4580267588269, 155.0107219615143, 154.93339049006002, 153.7810624077033, 149.54808846504, 157.19871468536635, 165.5289790518782, 172.3072755353122, 176.4788685690755, 184.27074797598794, 189.471062297489, 198.768566896243, 210.02364258663619, 220.7796788604067, 230.32264024374288, 236.90170679915968, 240.83312379139167, 247.79042677248862, 252.8989036208959, 257.59467652291056, 261.07363935732087, 262.80563589311447, 266.9465665915875, 263.3351927318172, 261.86783300522507, NaN, NaN, 29.00889033405146, 29.00513163173825, 30.472648941606057, 31.385574198453366, 32.59299960601854, 34.46302405582753, 35.30358700057145, 36.21971635898445, 36.50574512541664, 38.88572485681904, 40.01796397928425, 43.906597414722214, 46.94969883753348, 51.46111804798033, 50.681714442154316, 52.76369550795532, 55.43235291941152, 57.43782735680895, 59.33283180332092, 63.330057553648594, 67.57658355212297, 70.86661800212931, 74.27069467727554, 79.21815531719324, 84.82358095940383, 88.44503661360518, 91.07985160562933, 93.81995281496393, 99.42997126138363, 108.54549967329436, 109.18592304659876, 100.26763754123822, 97.07208875013309, 99.69952092430515, 105.06861086593216, 105.27970068288936, 104.28474426991424, 105.81588677607496, 111.31332741282148, 122.95301121284395, 139.2664833626958, 154.96078325937575, 157.87683934493583, 160.50819743022964, 160.52228198847666, 152.92867722213572, 148.13390493291766, 146.2828212494159, 147.47380431424006, 150.33192864908912, 157.2371731804497, 166.84034449412502, 173.99035330794553, 181.5516831471515, 189.79159795924343, 204.3772536839181, 213.94813242660652, 221.52062130743633, 232.38166279006865, 242.56981893563105, 249.02767667871677, 257.294826467995, 265.4060014129474, 268.6227268796744, 269.77230633437966, 271.01907108698117, 271.1386577390909, 270.0296527449007, 269.85433509804307, NaN, NaN, 28.891365624813904, 28.445686057869533, 29.472959745595155, 31.30755934723005, 33.73274993565434, 34.68239014067205, 35.41197442839707, 36.290151384484616, 37.23739323806076, 38.402699934712096, 44.200026423324225, 46.32277989186057, 46.53496309399756, 47.33458255044865, 48.87025847523532, 50.0334006911788, 52.22661826775417, 53.8327699216779, 54.48702788649903, 59.32548972190588, 65.22685959946689, 68.22610893489215, 70.34080794126962, 75.17576973966139, 79.05268311484593, 83.00392369340399, 85.48742417830047, 88.5574534731768, 91.84170623878002, 94.24919239923457, 99.07628683682341, 103.6083977659732, 105.1340082984013, 99.79515877450275, 95.9066413009588, 92.74762559176, 93.75281200411035, 97.48091204614565, 99.96322929443552, 103.04024496624291, 105.70134997302029, 113.18725031219448, 123.72319765897582, 135.8835327500452, 148.50123973206053, 154.79143841040448, 147.62190727859308, 151.00745812547726, 144.73176817801746, 145.19037624438675, 147.42723552412497, 147.78988409700648, 158.022736092824, 166.7569318346389, 175.3794166893356, 181.08911141149318, 196.2854661328335, 205.35785165767157, 214.72190157040632, 227.2379508405614, 235.81652250067995, 240.38513210978317, 252.26465680353138, 264.9591952160607, 266.76961410528594, 265.655858759098, 266.44742718776746, 267.8641576372075, 268.36745947516033, 268.42592965061556, 268.59693046478276, 268.6561526050751, NaN, NaN, 26.786906780007655, 27.078634561516242, 27.958809049789835, 29.279109098084028, 31.70044702995172, 33.53142693271196, 34.041690331985976, 34.47541700710648, 34.97902613199619, 35.70644879048074, 36.287481907126086, 38.043162583250165, 42.52002904203756, 45.81865074879534, 47.57273927644343, 49.398284728439194, 51.595725881999826, 51.58775914959697, 55.547103418801484, 60.826242394137786, 67.10006399705587, 73.03867349212777, 78.08577035098611, 81.30483472474972, 84.81833279869416, 87.0884103335547, 91.55662753838118, 96.97297964715642, 100.32960872761855, 97.25339586452239, 92.84990038667684, 93.35143683338092, 93.48606985617458, 94.35189849542928, 95.44557934283928, 98.4475166058699, 101.06619605133075, 103.988171141423, 105.3697672106468, 109.47014330667967, 122.47694263238539, 132.2942378539403, 145.34871873950902, 156.04852859213963, 148.01881382155455, 143.04265014626452, 148.19134624450814, 150.584146070588, 152.2707757873897, 154.5562471546707, 159.61018197154007, 170.3990690841975, 178.2016327842939, 193.3443826842057, 197.91315125477664, 202.92494224973777, 212.89922852576078, 222.98057633626732, 227.89669351804207, 234.41568432151502, 240.263365075359, 248.16827767435663, 257.0827895103337, 263.630552799151, 263.7338987695839, 264.3613581011897, 262.01603781852253, 259.3549068040143, 259.3850024078714, NaN, NaN, 27.639062807536494, 27.599004676865235, 29.02988880798789, 31.526707720386625, 33.03001010915282, 33.836240034533866, 34.126877385044466, 35.22422406964607, 37.79199451979346, 40.80182066230018, 44.105257198936314, 46.56132247862611, 48.28172924674167, 48.23698980610648, 47.16355530725776, 48.39829535622255, 51.657604948939664, 54.66230084750349, 55.49861445139444, 59.97214928621366, 66.27934578623571, 71.1143228569629, 75.80612050773976, 80.05376370162608, 84.45345672009441, 87.45289039042886, 92.0714670545912, 93.76137114152948, 89.94524561587612, 90.37366961240473, 92.55752054105527, 93.79559533967047, 92.16954171996574, 93.84098334474305, 96.9871275852635, 99.24454715389382, 103.26971927986756, 106.70416283908854, 111.08481735835788, 114.08651168200008, 124.17481984315873, 132.62647585706063, 141.1196247797489, 130.91554086773633, 135.42414783736413, 145.2531216766153, 149.4433488253551, 149.4765488910058, 148.4428599571035, 151.14276223440862, 159.22842900686408, 166.64158231426552, 171.79088877327487, 183.77282595828817, 190.93765592676053, 196.08032058819495, 209.69731768799008, 217.47237579167827, 223.88926548647376, 229.94879307934195, 232.39325843476158, 236.0696031734343, 240.9583143404874, 248.7273838441337, 256.7830539503586, 262.0875308198381, 263.0292560329714, 262.5779703580699, 261.5869632586885, 259.5366150024244, 259.1574318968218, 259.19260978671326, NaN, NaN, 28.52498671578619, 28.00517024745148, 29.25146690530223, 31.823483699875258, 32.92360375030312, 33.35657012105753, 33.9371383563518, 35.03572189757872, 38.631083573165185, 41.343046442044056, 43.17135078288088, 44.267038723809414, 46.75503709252851, 49.16842885244639, 49.45395933647136, 51.94347918830484, 54.65261994432812, 60.588110342286306, 64.98815108500351, 71.2222030363649, 73.78934394370569, 75.64849620735222, 80.81488532993617, 85.64417140125104, 89.82575432205327, 93.24507793936164, 98.84216911002395, 95.64840501780779, 94.09686037702492, 95.29809108438961, 96.39634908601604, 96.18561195442757, 100.13979119242329, 106.07426711852095, 105.85750243234546, 107.60637920850068, 111.3310748605443, 117.7012912222136, 125.05245030881692, 136.46542430851858, 152.22632512170605, 158.38093961891724, 152.255394052394, 141.47921885673375, 142.00199896065902, 148.9629960949979, 153.26047896691685, 151.2902781778024, 149.75691707860057, 151.74908118764296, 156.78267333696982, 164.32665711548185, 170.4918085749186, 181.27923485579103, 190.64787862882744, 197.75121750800415, 209.5123016402387, 222.63928932624512, 232.20118084378078, 239.92964194049722, 247.2551181385628, 250.82876446957383, 253.4715606785827, 263.4153664474755, 265.64826943601025, 266.21424312659445, 265.65021290806465, 263.4019842429638, 262.111001938787, NaN, NaN, 29.294961824789322, 29.329411141288514, 30.57707017091724, 31.195341024474757, 31.777921875824127, 32.581525976867816, 33.64113681003674, 36.428558373436765, 38.33294798230909, 40.45995245117904, 42.839541754631874, 45.84323312607649, 47.305591171504254, 48.14644854572948, 50.85733140310887, 53.08462411069388, 54.69294759851628, 57.02954089689667, 60.688364227948576, 64.9715702840759, 67.16693289821782, 71.23309221924201, 74.3075670969928, 78.59407199666337, 83.86609339030208, 88.48300982348775, 91.33107476423045, 86.05149162725917, 87.3674854847084, 91.86127239391256, 91.84887926594426, 92.50742580384563, 93.27653534790159, 94.92050989605329, 103.04273164254138, 108.75889319173046, 108.97932775762266, 112.15458218627177, 123.23998148675075, 135.87049708376327, 140.14711977825525, 141.14438047879102, 134.70672306716676, 134.7350148000045, 140.88028010078682, 144.8372720442501, 150.14704352161752, 150.91273639761062, 151.69882085062397, 151.18050120626273, 156.09102576694144, 164.50045381574517, 175.85480348221637, 189.24740855337134, 195.71638023094116, 206.01115320746783, 220.99408070516319, 231.83518539005934, 240.098058302954, 244.35130409589627, 246.85076794390295, 253.1454835047608, 262.18237771463504, 267.07126799055663, 265.357352668201, 263.10690167000604, 261.4987439587471, 261.4978843229556, NaN, NaN, 28.447703567893726, 28.443343679211637, 29.24723745428056, 29.90505944470763, 30.781433842395508, 32.10025406788232, 34.52082749604277, 35.7654320259669, 37.67178176919075, 40.31158722181904, 44.49685902416003, 47.35342911988314, 48.232963618849126, 48.6663738955988, 51.22693554114829, 53.425212980696664, 55.10284630763825, 58.762248469305725, 61.615051041416905, 66.67226933865166, 70.04532436687387, 70.91361361910866, 74.56858956772003, 76.90168398137669, 79.53666546193632, 83.78332239718833, 87.28698711189077, 90.50560081550111, 92.84550975698929, 96.35141796020132, 92.98073821811786, 88.28102298651991, 87.39187129740465, 89.58933082940202, 91.18789067693993, 93.08838746203845, 100.4286492045823, 105.84586413464879, 116.2626411294246, 132.53050312564082, 132.23625030723272, 127.85113546854694, 128.27419355307447, 136.62913325170842, 140.59522804919206, 148.10247353482777, 148.91500964720157, 145.43630162429298, 136.6841386265743, 151.27169167952283, 168.2717288613961, 183.302811610664, 192.84748267543122, 198.0587953400272, 209.3749369782718, 217.37066692471308, 227.7456728679839, 232.42118759972274, 239.4277705163468, 240.91921067186172, 243.38286289879755, 250.94436739393754, 255.86319100785406, 264.469342422195, 269.060538661127, 269.92152763653115, 270.00243538163465, 269.65486343965875, 269.63072317203944, NaN, NaN, 27.602363917459126, 28.114012993093386, 29.728958544703616, 30.607511742655774, 30.749851009355055, 31.111150428596254, 32.283829108267014, 33.60387868264241, 36.613256363861886, 37.85611302298136, 39.242385231918824, 42.467789582988985, 45.54609247007393, 47.670865088624836, 48.69238166784625, 50.73975260512672, 53.818245353730724, 59.61081830214427, 65.40396738665558, 68.69752907917041, 73.10314655935846, 75.47971663583768, 77.30433916106462, 81.33544322331072, 87.56014148492241, 92.15061005558522, 95.44593797289731, 91.60001526404875, 91.95745688848805, 94.50295231175922, 103.66053637914995, 98.52611088452518, 93.93360042099289, 93.91991979012248, 99.41452563998206, 103.80873064132572, 104.17659355285278, 115.72742034406056, 136.43729934167257, 140.26766612724785, 140.6392885423689, 149.66593903688386, 145.06811421447472, 144.6380337183529, 148.9423912589757, 148.30727042255953, 147.43997276818493, 145.16686005241408, 139.1416884103494, 151.61826391089005, 161.16852224831973, 172.91251228264525, 183.3691885812418, 196.5193589452171, 204.29871054957354, 211.01416362384518, 214.75536308432888, 223.02091322070729, 228.5064600152822, 232.66565464744988, 235.63869359839458, 243.32802117966216, 253.3584336769585, 260.5141545135277, 267.7575708767624, 270.67227381924715, 271.10901760617105, 271.28209630273216, 271.4671409765505, NaN, NaN, 30.892046886461305, 30.668514317768114, 31.76926158394497, 32.42345859775959, 32.85642866275736, 34.394217720470735, 37.1090236279318, 38.94044913631486, 40.47700224554626, 41.86527651212652, 45.83004668740319, 47.88055087349495, 48.31371983112434, 49.69979023017, 51.23568789727208, 53.06614119716689, 56.2910621773356, 60.466939868704515, 65.37774486962392, 70.21736879161543, 73.40123963068473, 76.80656576622182, 81.09469748056163, 85.16005893782062, 88.4486309683863, 91.62952836245344, 95.69338950652327, 99.20223875583986, 101.50587396343539, 98.53066625141625, 95.32515725126756, 94.97300453334609, 100.45812077125285, 98.68965398518502, 98.01561858501636, 98.22699374344876, 99.43568199195501, 104.04364694254366, 111.94359518375883, 121.49769722318217, 133.11658013745134, 143.39603639429572, 145.50409471996716, 150.78274870664092, 152.2326376819026, 150.6160090974326, 152.38034779081516, 154.47057023943898, 146.7545429423723, 151.8137893134011, 159.525460208, 169.02512458414085, 186.3664781189781, 195.04641610652374, 202.38764219978114, 207.07577924986234, 216.76206390599177, 225.48022546677257, 229.5912543541479, 238.78362695455476, 249.81782096202812, 260.34386214179165, 268.1833473690269, 269.25015678698173, 269.8396088881017, 270.5696890540816, 271.39534186683767, 271.4600056310923, NaN, NaN, 27.158764841618012, 27.377620524376713, 28.183406114785864, 29.430612872792945, 30.528078728658922, 31.996126928775166, 34.71259766510334, 37.503476104973295, 40.58751865312512, 43.44919542686688, 45.42624480604316, 47.405248063366365, 48.50434918563723, 49.96412124514909, 52.60044531912507, 55.16024187257815, 58.528870130840495, 63.95357814707122, 68.57380173264212, 70.9868111919025, 73.76599605794237, 76.62419331360077, 79.25968767009563, 82.44225421406317, 84.96341486383174, 90.58178446732416, 96.84194795149149, 99.9165442066455, 94.08202429330376, 90.11566325224148, 90.54593718046112, 92.73600090349771, 95.03674319989081, 98.42986967624843, 102.70674208035692, 105.33817143874505, 107.08530023436023, 109.82641460268627, 115.96555064338698, 128.0563246280276, 141.20161428519089, 154.0699458435382, 152.88377561037893, 145.48983785382484, 142.5232139918116, 144.82296504443997, 147.06777950830497, 148.47191573574875, 151.08031505662717, 154.08254989780164, 158.67592891901526, 170.66685275937746, 180.64983947737454, 193.35636417810744, 201.77987966453858, 207.29857961945405, 216.18259127391957, 223.68048570550354, 230.6853310279033, 244.47491351374865, 254.93152003447068, 263.9826198816795, 270.8418383600525, 272.6027192112787, 270.26007721248664, 268.4621840960995, 268.4456735113637, 268.52798103134927, 268.70873764334704, NaN, NaN, 27.67291951957633, 27.669720387800364, 28.91822918555626, 30.382250338488163, 31.554973260455796, 33.61291790852779, 36.84511369238473, 41.620116280395514, 45.14503275864608, 46.45595707545708, 47.772118740026436, 48.6443082759797, 49.73576175316118, 51.99925113063196, 54.560046952305946, 58.88152693104854, 61.58856752678709, 64.66057884865505, 66.26950533936258, 68.6112162751908, 74.8447243070883, 80.26275406225565, 85.2442545728862, 88.31890837610264, 92.8562045947322, 97.39208290913938, 101.93538215783516, 105.88217472433824, 110.56507921502067, 108.36788134641806, 100.1549486466924, 102.35756415777055, 105.72888546518156, 110.27106380840874, 114.94546234960575, 122.27075385730494, 133.40142566345642, 149.5276481162694, 146.75081446163108, 136.32699022841467, 138.43778915475943, 147.27526831938727, 140.98590105182163, 144.53085458296897, 150.55151090717413, 154.2405801112664, 159.57892595307527, 169.17444702050688, 169.0965125309406, 184.89683375865144, 195.7780045372054, 200.02232346906726, 206.5215445962156, 218.35796955637366, 224.68903430459292, 232.1301325894003, 244.2714247196498, 249.88123630369705, 254.707637069918, 262.5619639866619, 266.8880035627217, 268.0884216167099, 267.960672350832, 268.0405125578632, 267.9869393194112, 268.19235496718574, NaN, NaN, 28.192276964051228, 28.151098617217936, 28.697664717273735, 30.346970766297446, 31.702393163884796, 32.8000773610079, 34.19072629998627, 36.61145538656312, 38.956502904554, 41.37377050674775, 43.35351300998794, 46.54335627089461, 48.88982854649701, 51.82092505524034, 52.95092708877916, 53.858851742366696, 56.78904198255006, 58.24697440948281, 60.55053478077101, 63.409304936404304, 66.44913708556801, 69.2978167023649, 73.91193623844615, 75.80750480009927, 78.87524629372162, 83.26387912160666, 87.94929566225642, 90.13987832347375, 90.6356774517883, 92.7465020433785, 91.58039349354378, 95.23537189062662, 97.864476903144, 98.37771412074581, 95.44479766107764, 100.28891344173293, 102.92408331497462, 109.00370746655061, 114.12640569699465, 117.78014360629166, 126.59172940963428, 122.64868816935311, 128.82639266656756, 145.1365923686595, 146.15446363748467, 143.51462509706136, 144.70576925106602, 149.14941801364802, 136.8860836972063, 137.33930699752756, 150.8841853387541, 164.76726259487066, 177.8521240054167, 185.177654150747, 192.19009789656602, 198.17720638205378, 209.39221277115487, 219.05839119814084, 229.63147373432818, 237.21111655053227, 245.56238055435944, 253.34038455287043, 261.311868865419, 263.51065937341576, 263.6145982536934, 263.84604243120106, 263.07250821079583, 262.97341958869475, 263.28841760246166, 263.30567883032256, 263.72163923262775, NaN, NaN, 29.812680785387975, 29.07187579356713, 30.097460818007757, 31.488514960919314, 33.17637433490145, 35.156941162374395, 37.50470461294677, 41.1038529425357, 43.96425901035084, 45.94285786153943, 47.9929564155141, 49.822170087514856, 51.796581387050594, 53.18313685132778, 54.499288989932005, 55.81262241576855, 57.86271854617627, 60.937169049493214, 65.55309357287058, 69.06497455498007, 72.94728615723562, 79.00072079731193, 83.39219941539395, 86.31130609578894, 88.50175050099362, 91.24084538970071, 92.8801575653487, 93.59938756915369, 99.64863021800923, 97.08264287613788, 97.63367448509905, 96.34501243324011, 97.25424915937913, 102.20510663854036, 104.95129130789039, 104.94511814705378, 112.63440713512317, 132.42338520864013, 133.54605661229024, 125.48707433883689, 133.4149126355929, 145.40597898503958, 147.16367788653972, 146.9576391645238, 147.98140669830946, 149.66428203474067, 152.0345559721767, 159.65136052172107, 160.05472117282596, 166.63944212376651, 174.34757366253976, 183.22807070685155, 189.87369953768092, 197.52919162135802, 211.56121378945934, 220.40057249660373, 228.99305788023833, 234.71845106069952, 241.30889174319896, 246.57837438784023, 252.3855655796199, 257.02676435723174, 259.2967514502339, 260.32901419871894, 260.1069374301149, 260.6552117189936, 260.60797272990396, 260.170847412071, 259.4038114716938, 259.3274752466486, NaN, NaN, 31.33053580885449, 32.211089619798656, 33.45878947352373, 34.92554927663477, 37.49405848619424, 37.41271734687248, 39.244500635271876, 42.10753449886491, 45.41341172307818, 47.31708856628804, 48.853162917453844, 51.4892224132168, 53.53765175000207, 55.517970823951266, 56.766885189810814, 59.69142800599789, 62.54953264668127, 64.7405704170778, 68.47851836062232, 73.5379063532932, 78.37180219691744, 81.29868814225692, 84.07659590402295, 85.3794736870084, 88.30746005803022, 91.5324996272295, 97.40179425748686, 101.35995630300765, 103.41024855279376, 96.51180654831643, 94.8959846293778, 100.90517123480397, 103.53185167659632, 100.88282646366048, 99.55198950025984, 109.51938029383328, 127.8336227045113, 136.47798309637383, 125.48654256226591, 124.15614443967975, 127.96280916507575, 130.1805659530887, 136.76951612597182, 147.55651755778246, 150.84055157605633, 149.65115394996184, 148.12664044953556, 151.9005758696731, 152.60894965644027, 157.09599736473763, 164.56247908534704, 172.58892064667216, 183.7949962789258, 195.48040694908627, 207.08387437943546, 213.41864813515437, 220.57502300113464, 229.32047313814567, 236.40979897844818, 245.61169221603845, 252.9616974612519, 257.4600717561973, 265.3191034543224, 263.39318097775674, 260.39377378314816, 259.61517309657245, 258.81824209556936, 258.27466619039166, 258.4544674499016, NaN, NaN, 31.365182102832073, 31.914146500610947, 31.872592691672537, 33.40920107342302, 35.27941839666235, 36.44823010790233, 37.835793230126676, 40.218032377115534, 42.63522404924103, 44.57844076876699, 46.95721280551162, 49.52261707034607, 50.21327719851011, 50.82943425554702, 52.91524063551455, 56.87922777380227, 60.724012490906645, 64.6011430006482, 67.63710159889352, 70.41229291433906, 75.98032518603002, 78.61866581035943, 82.28637689694985, 87.85741406014367, 91.81893928100007, 100.03639820706498, 100.9158468618464, 97.53756063947272, 94.01095923706984, 97.09699092021847, 95.90114186721328, 97.78405758773062, 95.72051075112537, 101.71795012285533, 108.7373589055979, 112.40108689545723, 121.63450217292511, 115.62367399553038, 116.78668358077385, 133.35524130925452, 144.51274836103704, 150.25266346993752, 145.00194178071038, 148.57278086901144, 150.70948367816604, 149.99158518413418, 152.78656602902615, 160.47453242481285, 166.926289754113, 174.51556165514702, 184.82979867570597, 196.2834611590054, 205.96749937266827, 216.07576360098545, 226.32455143196927, 234.3079790332612, 244.2280349314749, 251.04405489315573, 256.75253093189457, 261.83658212423694, 264.63364777433674, 266.6670161293219, 260.85250774878847, 260.2198528818999, 260.75621848478676, 261.0237156500041, 260.52455393191747, 260.73140654117583, 260.8568479634549, NaN, NaN, 27.414628613217836, 27.30115887399087, 28.437641163824303, 30.384531438364068, 31.629761014078195, 32.72885528238613, 34.48839237243306, 36.175527901184616, 38.374659681735324, 40.49901731833262, 42.0010534987391, 43.5045242934321, 44.19574021289268, 45.108613990405885, 48.19056484595419, 49.874104386689126, 51.44616177694293, 54.6317438225655, 57.640397624141144, 60.609310569699225, 66.02853688302415, 70.49593510896135, 73.34935391512242, 77.23120594437592, 79.87114378993647, 82.79076780043897, 85.64563118296948, 90.33922899234754, 93.26768830491575, 100.23056266781964, 96.27085204261414, 91.05776191617213, 93.61279016867005, 97.99864666419923, 99.52297732132358, 94.30694074042987, 96.49693290753217, 104.26271872933414, 108.13779142940129, 109.81370683020205, 114.1295785292383, 123.21163645746104, 135.524708071858, 150.0424763616919, 154.60247242405876, 153.45225937976775, 148.65599965101876, 148.4167608307609, 150.06327066836528, 148.5246112398643, 153.76213607870363, 164.43968168248838, 174.2408670045854, 183.94109597435903, 194.39502160720463, 206.3484460486996, 216.0721291657789, 219.9785167846153, 224.41558561969686, 237.6339600429421, 244.30772982399688, 247.38693566384006, 252.08000022175978, 252.83660615074467, 257.27616906733124, 265.2973289408196, 263.73186255914305, 262.1100559021292, 260.7003650942101, 260.8105436657523, 260.859069473082, 260.9557795675198, 260.4176274699737, 259.54454093086025, NaN, NaN, 29.517491222163947, 29.955152990389735, 30.31895498581501, 31.564716557335966, 34.062681153329976, 34.79701132864636, 36.77791881615729, 36.846349686943945, 38.09068148080958, 40.73327242835831, 42.86126490508955, 45.57545339461457, 47.9968969590973, 50.26617824225196, 52.460431081859085, 54.79885375700322, 58.60942661426931, 61.322276757017164, 63.370502071531256, 68.12779291009979, 74.09931238205542, 77.61246985682948, 82.88661087425, 86.69394603534342, 88.29619212458472, 91.5146055679299, 93.85438036141521, 98.25088578360257, 101.03673856087346, 104.24853350943896, 110.54360212924549, 111.55616072725644, 107.31128766535433, 101.43983881321223, 104.07168998794327, 109.63492599648937, 110.0635438993963, 115.33082142597647, 121.34097047086324, 139.68355760526995, 141.92765629758722, 149.83268566151247, 151.82092714002033, 145.9418164805962, 145.90008751796438, 151.00272426735896, 152.2369957871402, 148.6795352561041, 153.97625106676327, 163.28899520126873, 170.40565324310833, 181.064876566567, 193.03074056543537, 205.3809305647291, 214.26367389453804, 220.79026289657997, 227.80099103824722, 233.12741568944398, 240.66716670669064, 247.89250194570778, 253.69457775427063, 255.4433634438803, 260.1904996317446, 267.1698332503863, 260.7509282226464, 258.443326443644, 259.2180347905688, 259.6194539068528, 259.94957806483706, 260.05897618599715, 259.39102241061215, NaN, NaN, 29.93113072225878, 29.411086540490828, 30.289475566829964, 31.093684872109932, 32.56034113063142, 33.95271768134722, 34.534174329856164, 35.04282139775605, 36.580094096722405, 38.85360180576768, 40.46840928218617, 40.75464852846178, 41.62998124882311, 43.24163658147378, 42.64880962096268, 44.1815686921874, 51.37934901828766, 54.16756835519318, 56.29481270214192, 58.05210987764547, 65.38971193681569, 73.15901713308936, 78.14341986549256, 83.71275345512333, 87.23403622674215, 95.14790128559933, 100.41493437089098, 104.80983392377063, 107.73371064527464, 110.07291776829572, 112.70823792562761, 117.0964828780284, 121.0447535745656, 124.26656728342238, 129.09489347734245, 134.6575663813855, 139.201427446759, 139.04909770997136, 122.0563961680997, 137.1704189884705, 150.5744879491982, 154.97867421283533, 158.39764917953394, 161.0304182093784, 159.5208743426925, 157.81857407078581, 161.75029142887473, 167.092841963282, 166.69858368504427, 168.42045008624032, 177.59610019102996, 191.2804702986578, 204.21195637203218, 212.32529713449364, 216.39813646020747, 220.87267529134914, 228.37874647890163, 235.23850977247426, 244.64688886067972, 249.94258168982572, 252.8771156270069, 257.36218439001016, 262.5060960282761, 265.3359315131765, 261.3786199839207, 258.7496880566661, 258.21359205878167, 257.84506880782214, 256.7413303110498, 253.9845476280595, 251.53616673420495, 251.28914327609198, NaN, NaN, 24.86011850466053, 24.707752097384418, 25.21719651844632, 26.535376726249115, 27.782579382348548, 28.36423268853234, 30.563846737537524, 33.28060201972819, 34.67110749721425, 35.47492179867392, 36.27992287491354, 37.89247542582037, 37.22926724780039, 39.06108784768996, 45.30576940273358, 50.59060338746174, 51.02644318890809, 54.69163695795614, 56.96522978029601, 59.16356828330819, 63.52677043402353, 68.80670739627517, 69.02082605258524, 69.7807561779707, 73.51840803319239, 75.60057549933471, 72.84479427135496, 75.36700636799164, 83.1737617315565, 91.96672779841256, 102.18950297325533, 106.25229800605935, 111.849413882956, 113.82652324024855, 115.91359496716298, 116.34505375874392, 123.37990518838006, 127.55152183513823, 135.0305395935658, 136.68055035752232, 143.6392329772799, 150.33533386318405, 150.66682784950996, 149.01017964871696, 156.40045704193088, 159.7344769123575, 161.41336853195165, 162.85243479288607, 151.3389596443726, 152.59396288125419, 159.78613999366397, 167.75628928519419, 170.37000828111496, 172.2563659866004, 179.0044595934592, 187.05104009432932, 196.16766935107526, 206.69781685275197, 217.12952461180026, 221.21827027683312, 228.16879753583007, 235.46838980730737, 241.68334438212784, 248.42750021817722, 253.23307930472726, 257.5741335134381, 263.3341927819941, 266.54329705750996, 265.1199593315436, 258.76612917415247, 250.87676697120202, 245.30571248201278, 244.5843226032827, 244.8364362165723, 245.24945767857892, 245.7331101866025, 245.91525588936463, NaN, NaN, 18.924304943659358, 18.99598382834656, 19.876851277775845, 20.82898642330741, 21.856284176608835, 23.178362686782297, 24.4235575429631, 26.69936039344706, 31.253830691639713, 34.41158283180821, 35.508294435393445, 35.72409956008601, 39.61858349165583, 43.732140528441334, 46.300923496818136, 52.171959654123874, 56.42192733474481, 58.466699358520415, 62.351341676027374, 66.82444697486567, 68.87144498404416, 72.05224494643498, 77.65949705237823, 80.51831270416994, 87.11211132435416, 88.98466293196296, 89.30996986384301, 95.36377837680642, 91.07328887978272, 88.63958809712729, 90.93512969039426, 97.086264426947, 106.00418701054437, 117.66181050394731, 129.86815838476423, 141.2139972671485, 145.0893027607916, 150.71905350261932, 155.45190735073277, 159.75535665618213, 162.44614819873206, 164.7967734752084, 167.5722314404933, 166.4161843665857, 160.20895588060114, 170.34223523737435, 183.25481009031162, 186.39276729626988, 192.09725824979705, 205.82391710954144, 216.58718701345123, 223.8715618368933, 228.12909549440514, 232.43979413947926, 236.5825963522482, 242.27551361617017, 247.69322387147824, 252.53022227192724, 257.4349966828897, 261.83530753450975, 265.0608308012917, 265.65971944669894, 260.8729722718502, 253.21934975724355, 246.40961721903858, 245.0430849982334, 245.2161468967253, 245.45980139902488, 245.55654349294764, 245.60152196399054, NaN, NaN, 20.87610049305881, 20.06223200844449, 20.794347596594278, 21.085632132157876, 22.186731848887174, 23.50942610702042, 24.53454305697843, 26.22278571770543, 28.349428785029378, 30.62427869655988, 33.48631999073609, 35.46694321737614, 37.59135363531703, 42.58376276796995, 44.93191578954586, 46.1751693930663, 47.417491523009666, 54.46593192939144, 60.19120684729412, 65.25174025364049, 68.07157071807178, 71.55249197048671, 71.90958595638809, 74.46972335534463, 76.1093795803053, 77.5715597881018, 82.87720604880555, 79.76212477243426, 78.28575157509867, 81.03318940164267, 86.53597750834506, 90.5616646158543, 95.1317187621558, 103.74134098370725, 126.09472827524189, 138.75836514442727, 142.60546052339066, 143.89796218712172, 149.3986652911042, 155.10527322957256, 157.65945040848896, 158.67547713926035, 160.93417585783635, 161.48367455375663, 164.36262032975412, 168.0463192083011, 170.05817317215119, 172.55516254896744, 177.59157620955162, 182.13357785068428, 189.83417981739512, 195.27716019340804, 202.70000270200802, 215.59675292244108, 221.87899255668358, 227.6284843170834, 231.54836132624433, 234.14438771785075, 238.66435046781262, 243.14505860054527, 249.3744218755969, 254.7576715278799, 257.8353763326428, 261.7678711070004, 262.88464168273754, 258.6108725719306, 252.70440364395196, 247.20173597492828, 245.8918947630398, 246.21612159973114, 246.38253522921607, 246.6305880742737, 246.80491738175988, NaN, NaN, 22.200442986649286, 21.68058091322899, 20.647240634326366, 20.936209852483696, 22.110359807445903, 23.35772336761646, 24.38432567717565, 25.1151791510419, 26.28788290035827, 27.679768990773358, 29.87903152796522, 33.10686563248271, 36.70524017142977, 38.90168165496432, 41.7621187010688, 43.51694573752623, 45.41909619702831, 49.087282245294325, 56.05962849534158, 63.845308202109614, 68.17869814244906, 67.407646841959, 70.4748208836399, 74.76328263710212, 70.57071439280817, 69.5665465735504, 81.00631615421526, 92.34218759143238, 101.91598005038307, 113.46999253419382, 125.24427051305805, 130.96348888842135, 132.15915469558539, 136.7886381896524, 141.06593837715684, 148.22975688835606, 156.612781648472, 161.45392257869858, 162.30918841919853, 161.41605989910244, 159.77586196218073, 159.1350376267004, 160.2731489153017, 164.26096526907133, 165.61489802363818, 169.17993831015002, 173.07443889360727, 178.15527906610257, 184.18243519065018, 191.0064140219342, 199.33083580817856, 210.9474131965763, 220.88555513723435, 226.46855714178494, 230.13873645704263, 233.77251513212877, 237.71059651500428, 242.50806471916937, 247.10007486924462, 251.41680175276414, 259.40392830359104, 264.3173873992593, 265.3153190297439, 260.86816063646444, 249.62209132198797, 246.15020194343307, 245.77470993655254, 245.76818823955617, 245.87658405756142, 246.18534462574112, 246.1509888383525, 246.22957145913972, NaN, NaN, 22.20084501606494, 21.901746469880724, 22.486540702410224, 23.438554581898945, 24.021020255573106, 25.928827389959146, 27.61497249276602, 26.655684753545955, 26.428750371318138, 28.629307887166032, 31.563984075786223, 34.86523622630044, 36.99497883827734, 39.93114743583165, 45.43840779144793, 47.63542816655024, 47.18640260441396, 53.64832335398427, 61.28714887136154, 68.78906891724081, 70.37081469458765, 73.89179032354228, 67.28172905935257, 64.40710160786881, 63.95601906501352, 67.13789886537049, 79.89919424265663, 90.46315022597733, 97.50153434855036, 108.93064984862293, 114.2075514904, 123.32407833995921, 130.80960094659244, 132.90522812699086, 127.17921088577246, 125.61972939704633, 128.14126874194955, 135.29281737479565, 130.3389271630606, 130.44818274944873, 137.42999493224892, 150.95747948184544, 154.0680581623295, 158.72907764357552, 165.02469753148665, 165.69436808772832, 168.68931106707072, 172.16857076832446, 175.5504605016619, 178.48023552824316, 181.76741133305737, 188.8032340804511, 199.3181634431779, 211.7150315729294, 222.7357641585806, 232.070131560677, 239.122460552318, 242.05093013240176, 248.36114404889523, 253.89554156090804, 259.1126938344167, 264.16379152837084, 265.3476012437674, 261.19740755745954, 257.8427806755656, 252.40038339909864, 248.06675314676215, 246.2362073513607, 246.0453302040677, 246.29741425851205, 246.4793011377712, 246.51506991903153, 246.6153499668828, 246.72377215305835, NaN, NaN, 23.166889186431472, 23.38431704072588, 24.484396595501746, 26.247086564455977, 26.61134014123552, 27.34455334553215, 28.445900355926852, 30.647154158512734, 33.36397275326049, 36.74475720435334, 40.12363711995456, 41.65915083984816, 42.536773218837254, 43.92237094467899, 46.48767483914957, 50.812966492065186, 54.335898516674604, 56.75271743508101, 59.61055560581119, 64.60572152848991, 67.72600995234461, 69.63570191434417, 67.72601447658202, 70.21833262298276, 73.44280013563764, 82.82626220172146, 84.13863117525192, 85.59108795423265, 89.25293189262493, 91.59368148775046, 100.09993921722693, 105.66992829670714, 106.10135419902103, 109.61346121130578, 114.30560465035525, 116.92589509779255, 120.00347705835426, 122.21569882491954, 139.96655057840073, 152.30510056299877, 148.25407776649413, 144.10352931595696, 147.79484091915452, 151.7215654001228, 157.97487982362654, 162.00246422547193, 167.8123853110545, 174.746979767474, 181.10091163461968, 191.0172895863629, 197.22711879975685, 205.86400600686056, 217.46073446974796, 229.31812805530592, 238.65004003116184, 243.39083894392456, 246.10199751592404, 250.81965888012763, 254.89163448737142, 258.906100325495, 261.6202051818217, 263.7656743017127, 264.85744887478313, 262.83872798565034, 251.50876777894987, 247.1467776550061, 246.8789726500243, 246.94707021846563, 246.9032573528872, 246.97957913728393, 247.1775325582342, 247.35748263475003, NaN, NaN, 21.09855399883189, 21.022499050380123, 21.755731643092886, 23.590507628115493, 25.206981265874223, 27.04271205149921, 28.584894532367542, 29.83275179287776, 34.09418211413629, 38.653418516980814, 40.70820937474256, 44.67058818581796, 46.057039623023336, 46.63509937941788, 50.37455141808926, 52.49331739893243, 54.614597415042276, 60.04413627288467, 62.02504944516385, 60.630850332242446, 65.8408010437809, 70.57371260924972, 70.56819474013226, 76.7320907338153, 86.53080152810739, 88.06745743748115, 88.49599280755099, 89.48392607504606, 98.49750876724153, 102.77748170995064, 104.43360963020677, 109.82176167027097, 113.11716233092241, 118.83262590709064, 122.13155458546031, 130.9375292832462, 138.2062343099236, 137.33227520460176, 134.2677889800727, 134.39940243667442, 136.44010115346302, 141.32022716574, 146.03554027397377, 153.47875195768574, 163.04654355765138, 169.15830140500037, 177.31730249352418, 182.2048875933999, 189.73295377471527, 195.65683893087066, 202.5271038282884, 213.3526944020988, 225.6533443873151, 233.53845608289382, 239.255401141471, 243.629155408868, 246.88032119290975, 253.42130431721503, 261.1052971398116, 264.7327367191347, 265.6423403806373, 265.09638826170914, 259.83527497802714, 248.5785176437958, 246.4185343493119, 246.3657573403984, 246.65171836615855, 246.826759437204, 247.1144167244382, 247.085340426097, NaN, NaN, 22.981929646030984, 22.75830167298224, 23.712731909150023, 24.963514379218495, 27.243342312489315, 28.269057359799163, 29.145898412554622, 31.495564123804574, 37.23262713080162, 40.02700102745236, 40.38953976188511, 43.83940515615798, 45.74364833562721, 46.98500083872521, 48.0761825681374, 48.72561321117473, 51.513230244347355, 53.9292538436788, 53.778797200070606, 55.67906371809176, 61.39904067277811, 67.99739682801011, 68.97990001155307, 70.29284148403433, 74.02787315659575, 81.61058938858528, 86.1143163583216, 88.5251655771725, 95.01793944159718, 96.67036321673397, 100.19103550313085, 98.87012220027958, 101.06543368043673, 110.42865792069523, 116.38257833978041, 120.90915369194113, 118.15019494157252, 117.70263547032732, 121.12309073874763, 116.94296304917901, 122.45081648796645, 129.84920352984608, 134.1662425587323, 140.5701547200059, 146.21880201654747, 155.08791447813434, 162.53364818329058, 171.34454305767534, 181.30734627307004, 192.29237633354774, 202.631609230588, 213.03488641946402, 224.87152909404608, 233.9700103853205, 239.24176198351103, 244.05958306645516, 251.34655353641915, 257.6489533105248, 262.3119218691497, 264.85043731041713, 264.327608292151, 260.9681342166292, 249.16259842111364, 246.35347292745232, 246.4126200814761, 246.6879607333546, 246.97867928241695, 247.25909298900766, 247.32859716060275, 247.4168962021368, NaN, NaN, 23.462550647800985, 22.79821927741868, 24.63770958783008, 25.81343699652533, 28.240051294846303, 30.960136705563205, 36.401370866636455, 41.846519994615804, 44.04919252144547, 43.89470773352213, 43.44506751667931, 44.61220807117898, 47.83988143137432, 50.84427927673305, 54.065779179439964, 54.71971419344998, 59.048129556045794, 59.99624856320757, 63.080083131704285, 64.61965029417723, 65.75042604878934, 68.05764734981683, 68.60214395649554, 69.14551191843438, 70.0214170907575, 81.02826892140921, 88.29132972959597, 84.32733025384108, 84.87297220638918, 94.33183314720041, 97.96908170634056, 96.7531558745725, 96.31126544401545, 102.5811985836441, 97.07064669092759, 95.40830964666016, 92.88073381968658, 98.51269862182278, 103.03256020484278, 107.98429788400577, 114.14621673657226, 122.29830773855429, 129.2510969963656, 133.00673908827315, 136.43098109224118, 139.7347439874262, 143.61559788484112, 153.17714891993924, 165.2787244146202, 174.52384348691044, 186.1781515508955, 194.00199102223283, 201.6644362255069, 212.82388032036135, 221.19086015987992, 229.54774949035044, 235.0396035366282, 241.90449530644864, 246.61795383135984, 253.31672644166017, 258.1038691062879, 261.7405824442101, 264.4202761670562, 265.63031675808713, 257.2973385318339, 247.04039865809307, 246.31229308201284, 246.5953796670776, 246.8906136434764, 247.18114660502434, 247.24193703826685, 247.4142050878587, 247.49779550280007, NaN, NaN, 22.505213602148796, 22.42889666993244, 22.942522290094118, 23.75004987696561, 26.76340256526097, 29.11413878810644, 30.72721748995113, 32.48893202501309, 36.38375935706396, 41.379244678234336, 44.025512959985846, 42.03607670757152, 46.07299683873601, 51.65389785846591, 53.92437363005578, 57.95282714382851, 62.19864498088045, 63.809571976338106, 64.46797660346233, 66.00983677137556, 67.24815765038188, 68.34304552091069, 67.38423391738948, 67.81668513723443, 70.7447856373265, 74.3299842828641, 78.4369802281599, 80.93187445335064, 83.79427733964431, 82.69127496723328, 84.0743413564585, 82.22960309231078, 84.7910696520844, 88.23353170354999, 92.12580292502398, 93.3713026575274, 93.94820583695999, 97.02647826063097, 101.14590861122308, 107.55251949124258, 113.8006843920623, 121.64320565845121, 133.0000226329254, 138.63742705612393, 140.53791267961302, 149.71858504171183, 158.17316458935457, 171.3148046779796, 185.30696303530937, 197.40573586545082, 206.20268636661407, 215.60743094950902, 226.65941922771793, 235.11966847201185, 241.3399804487701, 244.12245208941388, 248.93506749916165, 252.83625725556598, 259.1662334819858, 262.5732296948567, 263.92456839004336, 265.1916678149622, 259.5624763606167, 250.86469938394066, 246.00980644608907, 245.52191257910664, 245.70406803728673, 245.8777620303064, 246.13535679389383, 246.2428027169555, 246.27480892453818, NaN, NaN, 22.541847962427823, 22.833841528944227, 23.787137818299716, 25.62281146703003, 27.533437603689368, 29.148141544411324, 30.246269034290762, 33.332362540355625, 39.21042471778826, 42.51548094930167, 45.819312670782274, 45.37663276928218, 46.17838844521669, 48.815810464065386, 55.27723249980378, 60.85778323725934, 64.08333730298375, 66.20972358641744, 67.0097104080823, 66.41351030071283, 68.13303936035646, 68.35018246747686, 67.17213025569878, 69.07265053325258, 73.02883911154962, 77.35823948949516, 79.92228823063614, 80.05836411243276, 80.56513745180311, 81.66295764988485, 81.59051201470928, 83.0530277464673, 86.27262253144406, 90.45126408841519, 93.01331869076823, 93.73755416425978, 95.26764663525006, 97.91459746043378, 104.46030777905831, 111.90401251520201, 123.9411215996895, 135.45865027252503, 142.13573214593254, 150.7593679365932, 159.1786360649833, 167.22389009350604, 178.70735826397203, 188.68889018737963, 199.02041514993638, 206.63629635370842, 214.22326560526184, 220.56645786998607, 229.55473653646962, 237.61909310184703, 242.79125600631545, 247.73336763836485, 253.16791787390656, 257.6813959818153, 262.74379158130165, 263.0753776717381, 257.62141857031287, 246.8753620552539, 244.62807332072703, 244.9154661471154, 245.0926568846829, 245.16157106369045, 245.44480003422663, 245.39103748439516, 245.33686523396563, 245.39804011180365, 245.36699809648258, NaN, NaN, 20.254207966654533, 20.39874216839722, 22.23761005972271, 24.149602634153254, 25.027946563639144, 27.231534317260277, 28.330682069577374, 31.48948676023735, 34.86834344989112, 36.77274739758477, 39.56349409757586, 41.1769552098004, 40.36572695731832, 38.96695955436692, 38.00820076150889, 40.64869269843239, 43.876571315971574, 46.293763820530934, 49.52050708057159, 54.66243455989587, 61.634080499641605, 66.62220908333931, 68.30872894962461, 68.08449176251635, 71.46430866869368, 75.20871724060262, 74.5426615942369, 76.81007846308202, 77.75776661492975, 76.72299458600419, 78.62646958472969, 80.46343212939631, 83.24635471404429, 87.13137488515837, 90.5060730406549, 93.21311979678002, 94.75286402459389, 100.1005908350484, 103.46468385387432, 106.18410832493073, 111.88509091558504, 114.55177262723011, 125.59089615148885, 134.42525844135284, 140.06512075833925, 144.0649194708739, 151.26063535090367, 162.16365338334018, 174.517087218028, 183.1005463430258, 190.25293184280994, 200.28183299752158, 210.47522599945353, 220.10809921116567, 232.53585808729497, 239.27204924590595, 245.59951063659906, 251.31967314975432, 254.30450164934052, 257.0116072286389, 261.6765344734774, 264.7843784305448, 263.7577273995908, 251.9251149882917, 245.77116086008414, 245.4973378270227, 245.78684677772898, 245.9551317024721, 246.12865660618803, 246.19876966377805, 246.37156013806066, NaN, NaN, 21.506913547434415, 21.393459985158866, 22.753254078178557, 24.957261818390716, 25.063053774668834, 26.05121379167905, 28.106270849025606, 30.41784632052852, 31.22337403257412, 32.87452449797455, 33.23968777941313, 33.16432114835062, 34.41360836782355, 37.9409187581932, 40.807774132877775, 43.96627650303876, 46.35100360241988, 48.258338431461524, 49.83345921480779, 50.746722960362774, 54.71503249726536, 58.23802171396653, 60.98736118254415, 64.61406178359029, 65.93288759517866, 68.67925745439274, 69.22682427727229, 71.7566581034604, 74.0587768499292, 79.11801230945315, 83.30584855662877, 86.27894649785885, 88.1434040235424, 93.64753349842977, 104.9739615843702, 106.50612046052605, 110.57257964990683, 109.24743296855851, 111.67625186751825, 112.00575492372606, 116.56532994306629, 125.83807986725782, 131.58455530571226, 135.90425833428247, 146.02792079902102, 157.03251792141427, 168.06737124758416, 177.96275160989094, 186.82023516457022, 196.9283982682095, 207.08389471711476, 214.26019010849376, 220.07977234637167, 226.14171370088727, 234.63021870996445, 239.3262447143653, 245.25231700893087, 248.1429010534356, 250.9071580256688, 254.33082055784567, 257.9505672926459, 263.2064038878629, 264.91515558088054, 260.21789321039023, 246.8558674823323, 244.1236043985401, 244.30883626691852, 244.70765583231758, 244.9929854006937, 245.06135012276908, 245.13317443983777, 245.32438945395674, 245.29084490136418, NaN, NaN, 22.509728710856734, 23.021563231555273, 23.975645431157645, 24.41114246785387, 25.363887219698896, 26.390693018260038, 27.41649686929866, 28.368884846171486, 29.430743666449033, 31.267494554113, 33.13666904444017, 34.674689198243804, 37.46536599262806, 40.99199203280439, 43.08241107747681, 44.284361711108566, 44.8276000421714, 45.997648835235545, 46.32185184379376, 50.21061742116222, 55.31893553311907, 59.17201230800158, 60.81701937357866, 63.34543884165589, 68.19507227984184, 70.93978106843123, 70.48870078246829, 71.91416434290565, 75.87941821382877, 81.93231140802914, 86.11050653544035, 88.96580430489745, 98.63761909472798, 105.45204307059254, 106.99192692874139, 109.73711518333518, 109.29756001224962, 108.96089863079254, 110.30957821821815, 115.81419196651989, 123.05463064093325, 128.02295485888112, 136.56529767077205, 145.11485982350436, 153.24185528826385, 164.57856852746227, 174.1345343735507, 179.79169683381085, 185.58546445121044, 194.69212470840262, 205.61996889811272, 215.69290994841336, 221.47248359654475, 225.0987129283781, 234.9203967364823, 243.0684757405874, 247.9325127606775, 250.89448790117177, 256.4534542671738, 261.5704940140553, 264.8406482716705, 256.84680249396433, 246.19896732653882, 245.24697658084932, 245.42453816920954, 245.829229073573, 246.0119266629656, 246.19300511887502, 246.24460145025915, 246.31732518653615, NaN, NaN, 23.35933854078289, 23.39323797170358, 23.684334851861106, 24.638572214017106, 25.740153727289137, 27.318614967184562, 28.674964889330077, 29.84724883073753, 30.721559576102837, 32.04050576280703, 34.79772710077048, 37.11113011974763, 38.650738922494654, 41.3705511722624, 42.320135551465924, 41.8702013002362, 43.59305086214687, 46.19604015204086, 49.49896398883804, 52.029322392050574, 56.8370590713831, 59.14837971233923, 60.897313043021285, 63.42317823643338, 66.51075707368953, 68.4892115710754, 70.35522538897862, 74.9853129733204, 80.49173610393505, 83.89473957250235, 85.75640871089146, 88.94780110147221, 100.2909524993053, 101.50282756261139, 99.51276101132575, 98.74607240666467, 102.71214522807108, 110.85784634971466, 111.86190345213839, 113.30724462622301, 122.67792289384529, 131.9429262498753, 138.47398060991614, 142.9262310880727, 151.92393843572367, 161.91686073825161, 170.47834917729793, 178.4731891306951, 188.94063743109575, 202.43168827659278, 214.04474802109814, 221.07223999817805, 229.70284322786767, 240.6531115053318, 247.32221661382792, 249.5648201525426, 254.29774303136807, 259.5719808318389, 262.31713949654943, 265.5352377735067, 263.2135264953792, 256.908200020059, 246.12081090579665, 244.712996356439, 244.8831644120675, 245.054308761606, 245.3433842040386, 245.4068157928042, 245.5912662428878, 245.66106742459448, NaN, NaN, 22.179641277196385, 22.2134251856727, 22.614693673204243, 23.123296291023188, 24.297146698794577, 25.95057355292641, 27.307597197720384, 28.516123508455248, 29.83636261844073, 30.862237429154742, 32.9169954153628, 36.14852007715523, 36.474926481143, 37.314749104415505, 38.63286897179388, 39.6914177511241, 39.75753942303297, 41.25552131246141, 43.527860691855956, 45.3626203122588, 47.5250731710113, 49.503869805796924, 54.45304675999722, 59.18449017147951, 59.72900338712704, 63.13768844858695, 64.67244881994087, 66.20940795662801, 67.8615115024052, 72.48635249127823, 77.33155439937158, 80.74252471137984, 84.3752260988536, 87.12432265937629, 90.8649091346338, 101.2058119927454, 105.27832298307369, 99.65938361848082, 96.78767391058858, 99.97226429422976, 108.41831708078556, 112.94138956984303, 119.9257323815951, 128.65661962417758, 138.8140588167478, 146.57297630047114, 154.37956823858337, 163.01805208586597, 172.50455739338588, 182.5627568103477, 195.14401833162435, 206.4203766826082, 218.80302417078468, 226.61317964793514, 235.3629424214423, 241.2746888664293, 246.4304995985651, 251.95838660446026, 256.6668225051575, 259.7029435303955, 263.2817463471218, 265.8029584508886, 264.9703022865869, 257.4292849218328, 247.7251836784315, 246.13041888541858, 246.21244379817128, 246.50567885842477, 246.58515415726382, 246.76817129913988, 246.8490757426858, 246.803281656632, 246.9845906350011, 247.05393516128575, NaN, NaN, 22.06980435453435, 22.25069831625517, 22.54283398497632, 23.82843836108939, 25.113602930606366, 26.250495272485495, 27.68269967782795, 28.743711143728728, 30.02754208001972, 32.305587883297505, 33.589709496816766, 36.01212579942271, 37.848270879889746, 37.29080744822159, 38.461652918031845, 40.036828256544446, 41.723545477436616, 43.664100358200805, 46.85394051031218, 48.5382129743265, 54.00042041367103, 57.44770728824501, 60.087015212227, 65.07817845515302, 67.87006450774444, 69.76968804517759, 69.40278579070139, 72.11250470206897, 73.58144022952261, 73.49901848957305, 75.54915762397215, 80.53363640244481, 82.87733434472185, 90.87960014497645, 90.87978835628576, 93.44453434491247, 95.93731248868494, 101.5972346247647, 105.48467773330083, 110.11283190488393, 114.30324496591406, 122.46537591076675, 129.63567510408637, 135.04586602615396, 143.3823248340356, 151.82743327038497, 159.80151424474067, 165.9372511437676, 174.61863100012206, 188.21447687946588, 198.35756280212436, 205.7010765516374, 212.88807502422242, 220.51163273789555, 228.4706621111657, 238.75170454740504, 245.50251826939174, 251.76132798656147, 257.00335163798076, 262.1036237325363, 265.44255686520086, 255.23597950482406, 246.1146562512004, 245.51548546374062, 245.69325752521374, 245.8673496368627, 246.14995365661824, 246.1087872148121, 246.18231182737736, 246.23837850889865, 246.29970097402122, NaN, NaN, 21.552086876000928, 21.216673611759784, 21.949647326774084, 22.68102696858928, 24.223402354520417, 25.581941671539976, 26.903331808256137, 28.33407007660837, 29.61766732239814, 29.979554508422137, 33.17455731594964, 35.92932378534965, 38.38694537231648, 39.01061613280909, 38.746620528903534, 41.35185522198454, 45.3509451446059, 47.76764407036419, 50.51860711381815, 53.45400723142122, 56.017222792712076, 60.425982072220776, 61.629526492873104, 61.73179427432842, 61.61621173682029, 62.15942034692235, 66.45197770066427, 69.09279333015184, 72.39247648721226, 75.35287386979776, 77.77173918768766, 81.5105964799315, 82.937842241206, 87.11927513457353, 91.52416129406535, 95.81347788731107, 99.77059836537687, 109.47562418712837, 116.10727005459421, 119.85155943730987, 125.88834456911661, 130.95833443961283, 136.1641277739623, 142.93150036631832, 150.58708395285666, 156.77706316247122, 162.769005642146, 170.68800545176182, 179.7031636804608, 185.60475955338597, 191.60595583348666, 199.43590975906437, 205.89041341899662, 215.4152774646048, 225.36362194711364, 231.87564427253972, 239.78301006919727, 248.19830591328582, 256.4206913980914, 262.566029065852, 264.65998552830064, 250.67381674623334, 245.20508092640466, 245.15942538904767, 245.56775270593818, 245.82079903971533, 246.0553151807456, 246.1565747537454, 246.26152598296883, 246.39582729735724, 246.35203461434247, 246.44835935219228, NaN, NaN, 21.51743195926257, 21.58692896538887, 22.54197836165633, 23.64151525083307, 24.962331608964295, 26.358644551837354, 27.017169623399948, 27.380445479727467, 28.406995592932933, 29.726905904149962, 31.55969659925269, 34.05530862370931, 37.873586372836066, 43.308576190709665, 42.42656109535647, 41.833299328006404, 46.6788964582859, 49.61077168810076, 50.560348824814405, 53.2683208657098, 57.051826242170186, 60.690446894581804, 64.43054583391996, 66.84723160623501, 67.3914749366788, 68.92976031544521, 68.81838548241795, 70.6816503740136, 73.98490027834411, 76.30012015718408, 78.05674377267582, 79.71400476317876, 83.45954078216015, 87.85307483499294, 92.69403730475318, 95.33441690577622, 100.28598702364464, 109.53850522856364, 110.09905290955578, 113.29536581056, 119.43988074246772, 126.833276154075, 132.01671115441957, 136.55015238882288, 144.21128974066744, 153.54671349580588, 161.97850868867715, 169.10152313424675, 177.92647314807428, 186.6460371515656, 193.9870642564888, 199.0713147660899, 209.4375618599797, 217.44284995181087, 222.27592033456233, 228.89810578975366, 236.25569005058028, 242.9997943070109, 248.5998800628443, 253.34858028274866, 259.4613952595325, 263.4670743334116, 265.80440418547664, 263.833901209962, 248.26368487629293, 245.21699185582887, 245.45781614716827, 245.70345491667914, 245.95582055386961, 246.20085052403093, 246.1449210024621, 246.2416746485226, NaN, NaN, 22.181154273646435, 22.177745556377538, 22.986480313750768, 24.45554544680494, 25.334077176823637, 26.068244546791284, 27.170425122153812, 27.829200027104662, 29.66645554013717, 33.928909998130244, 39.29444245755312, 38.70489537363045, 38.33020193557607, 40.01549690832984, 40.232563965199176, 44.78887731536421, 49.34568169768998, 52.05685701430277, 54.83956272856603, 58.21086291787938, 60.33380894484914, 62.82217460014754, 64.87421722898063, 66.41794830406674, 68.0342981006455, 69.35245926258725, 72.42763330581151, 73.74038489011139, 75.34879690378973, 76.96412704415195, 78.0624038786674, 82.39267151683318, 86.42966325636336, 89.86762527417993, 93.24037463482776, 97.1992412917796, 104.46092090706104, 111.43010612881615, 114.08632367126425, 119.26106643292754, 122.65851179674728, 132.51406420654166, 140.31685996448883, 147.40369428839895, 153.3166845458119, 161.47269695727363, 172.18131751642616, 179.72759452668325, 182.48663302155938, 190.24673441715962, 206.3213187061851, 218.89772601986797, 225.48547382286554, 235.38913582791042, 241.86409268103162, 247.67877342007955, 253.16651820747668, 258.12377978513456, 262.5790808561133, 266.0853272124063, 267.49456995410463, 255.39184952211613, 246.02659042125111, 245.5219603148008, 245.80765967158996, 246.09209563674122, 246.38364408721938, 246.44345674076138, 246.50747202798803, 246.45907224453626, 246.64869350839072, NaN, NaN, 22.659574609241506, 22.43503251540612, 23.574859919648045, 24.565595038832832, 25.484980513282828, 26.07038191950349, 26.8395973274023, 28.527486222023665, 31.90978828905038, 35.105421443972965, 38.08017363498967, 41.019028490395165, 42.04765909651955, 39.61718840906731, 42.26000784458895, 46.115487424929015, 47.618009793343, 50.59152355584732, 52.09228975425398, 54.44044406900788, 57.523120632728244, 60.23547799403534, 63.16695350497456, 65.14188596457102, 69.02987786575717, 71.44831584699281, 73.57580996724568, 74.66722689479664, 74.582351400771, 76.63427563047205, 79.49102536436794, 81.68902073544311, 85.79653313630389, 87.3225701697454, 90.558271840639, 93.11992875633547, 96.05989664323798, 101.12861834186268, 104.00297829425395, 108.11559615873784, 116.13378463915673, 120.9938110218438, 127.3344180297015, 128.40028279325742, 131.3611357214184, 144.93014170019612, 152.628249467362, 160.08332114545001, 165.33970198806284, 171.57592135555802, 187.58105033009988, 200.42603421387187, 211.36221545933012, 220.35645491756995, 224.19288618021102, 229.04421641729118, 236.44417673404354, 243.4641037675635, 248.09013547373328, 253.4604337705384, 260.06869523699885, 265.68175645741155, 262.9647087367898, 247.41546622447595, 244.8163651222833, 245.06945973387406, 245.33533618766043, 245.74447154203156, 245.85472702525567, 245.95809141309013, 246.06369812562664, 246.15859914015957, 246.2671574692858, NaN, NaN, 31.914327023618316, 23.651058605461433, 23.42674602251999, 24.30618198570963, 24.37740326934597, 25.55126002241868, 26.945839370381602, 27.453379572722106, 28.77253956670899, 33.6213145791653, 36.77752515621535, 36.55319776808464, 37.43265097528807, 39.852612895237215, 41.53807989315229, 43.22374278773691, 45.57044614011333, 48.13847365329119, 50.40966352478666, 54.446996951238276, 58.11446729999857, 62.59377782578855, 66.48416063767618, 69.19430276071253, 71.53462749824133, 72.11993380173521, 73.73209673527316, 77.39668636673606, 81.06953634431412, 82.60351273085891, 85.60970148856542, 85.75315367838584, 85.89983847759665, 88.90216830233975, 96.31783078365186, 102.03464258067035, 106.51264203702294, 108.4368778985816, 105.94795637636801, 109.75976406201062, 111.93644308983066, 120.9250331634437, 137.99612434564935, 146.4294860690064, 151.73586411075334, 150.45325973979547, 163.73235021807892, 177.29236417545206, 186.8355322487639, 196.2510906050104, 210.51061261902416, 221.1691137173806, 228.07031860678384, 236.06058077390884, 241.3342203552858, 246.61225941439017, 253.69237258487397, 260.5469222319998, 264.4808418040453, 265.6520115735831, 260.01169311206803, 246.03692960806615, 244.6364880083599, 245.04154281941913, 245.29769011369856, 245.55359697268378, 245.6695305104219, 245.77631085765609, 245.88110905080617, 245.9946466864515, NaN, NaN, 21.107047854381406, 20.88242928736921, 21.763713536215057, 23.233973230242338, 24.03952379523021, 24.439529524566716, 24.805178610163924, 25.610299441484607, 27.188461337311985, 28.72632574339886, 31.03796373759295, 34.78547965708568, 37.17381692169403, 37.83068320571317, 38.67085581604578, 38.95736240118404, 41.0090700421546, 44.31084831427834, 46.84387949537826, 48.56211207474978, 50.64904823865747, 52.920024719918736, 55.11791802141965, 57.39112833715409, 59.588608315528695, 62.66349284424034, 65.96489910059793, 69.85338174490133, 72.63912771385576, 76.37291898683456, 78.27796103996918, 79.59616915474056, 80.54850798086717, 81.13421423739429, 81.87249865417243, 84.07088382054067, 86.7836398086212, 92.13987042586476, 99.1893098368175, 105.5770006001091, 109.44123488240467, 112.76106215963236, 113.50714944325412, 117.57633478837462, 124.97599684854524, 129.9773714770813, 134.4281424014058, 141.80966572062, 150.11550204950876, 159.0131913922672, 172.03477115482247, 190.5427619074078, 209.8410088232296, 222.42252931212096, 232.58417465389354, 241.00561473786587, 250.13655124648346, 255.25389058106825, 257.9176912940806, 261.40208590830093, 264.6686932192123, 263.03383374521036, 250.08489310142966, 244.6087141067817, 244.67410477656014, 244.97231058556164, 245.26738634053598, 245.44975540727324, 245.62446295007248, 245.7990916078721, 245.860913154715, 245.92593241741193, 246.00726554774894, NaN, NaN, 22.989477766648317, 22.94924223846468, 23.31303269058897, 23.897943388308015, 24.4818408856641, 24.736854919926593, 26.537456668922985, 29.475135929794828, 30.724070083592547, 32.52082344483691, 33.76533539755377, 33.50496371881647, 35.00369811769043, 35.55229735237532, 37.42076759823196, 40.391233410257925, 42.588875306530745, 44.82343415064281, 46.80375396127157, 49.186747884112435, 51.16678516240718, 53.77182031809205, 57.76987438585608, 60.52501802271811, 62.321390047467325, 64.99506455102929, 68.40518267306223, 71.96187840567097, 75.36928547330366, 78.37679419967448, 77.38426882093677, 78.66904963603102, 81.09366369029455, 83.54273994868423, 84.9711721567151, 89.44870014990512, 93.40590407985191, 95.71752270110036, 99.94333938996085, 103.43385967755387, 108.13195531566295, 111.09160980175426, 114.79451574294258, 119.6724980406532, 125.58397658523718, 128.11329729840256, 134.47745186055943, 142.00566431822307, 149.28157513333312, 160.56039309813983, 177.85087896162784, 195.1338016265379, 208.29331149748566, 219.10482219514336, 231.28651143918307, 239.62034592439238, 247.74353938301164, 252.58553133863072, 255.68669241381807, 259.6147673927636, 263.65665582324084, 263.13398750613516, 262.87892823608615, 256.0246843086524, 245.4085281510744, 244.7908736627373, 245.08373306817572, 245.4848974976415, 245.76702765608033, 245.83954002094066, 245.90819855379812, 246.08668816824976, 246.0503684297106, NaN, NaN, 22.62274157353926, 22.619235238386434, 23.612879328467198, 24.418302127912227, 24.673898601011576, 25.479606551002096, 27.795337918359095, 30.73320810970917, 32.495728715759654, 32.89439540481508, 32.74307388558989, 33.65671625213185, 35.0854948943387, 36.366127077365434, 38.197651785155074, 41.577009379142055, 44.65885519124581, 46.3774811567675, 48.57646947954919, 51.7354633783102, 55.663506674071854, 59.921558728564214, 59.62890793210559, 62.04598678200808, 64.76109509554425, 67.10625195658463, 69.52158568259313, 72.81997884068252, 76.41071178884559, 78.68687075997755, 78.9817492729185, 81.02971126726653, 83.078926576732, 81.53651370250059, 83.73242172707893, 86.95934432694918, 94.38235854242295, 95.850456710784, 98.19612670656753, 103.42557502255217, 109.28920293221407, 113.56644182132109, 115.49403387510499, 121.41219366318705, 126.46273310198525, 132.3855584998209, 142.15608644190735, 151.66039088844147, 162.64661766364156, 173.19876806319834, 185.39491722067947, 196.7194658947014, 211.04905723645413, 224.96788596381307, 232.37824501085325, 237.82541899192992, 242.57825269154495, 248.53927713614112, 252.38888203480633, 257.15515571130663, 261.56907126463324, 264.75862729402303, 265.2723300565423, 264.70207284744924, 261.8283903470557, 249.9929903024463, 245.0772390999092, 245.18326441068095, 245.58533609910683, 245.76399486638408, 245.9431490683519, 246.123375294657, 246.0902800203776, 245.95883794151186, NaN, NaN, 23.989988878013605, 23.617581954890476, 24.203910985166328, 25.30613249822487, 26.408510762863116, 27.508886324818388, 31.479603090569018, 34.71631786849485, 36.405409122152825, 35.88603015668385, 36.470347200640504, 38.15701975308613, 41.609910551849595, 45.507563754877665, 47.55827277327393, 49.31554242758338, 52.104570610186194, 54.746275920928646, 60.03321605754302, 62.306433010750354, 61.644499341182296, 64.06597539776583, 66.25950311398049, 70.07861920842468, 73.45758888152194, 76.31581074207497, 80.20647099834665, 79.09858905116624, 78.6516811044656, 81.2168066497593, 84.66481914209112, 86.8612173882293, 88.47244015383215, 93.68025166901775, 98.2350356984093, 102.56680400040531, 104.91920857762176, 107.04313170536486, 110.5802941712832, 112.88080922760268, 116.56482770216688, 120.55947091988308, 122.66932404436253, 131.54721039701303, 145.0202679373003, 153.0439495964105, 160.9001899357502, 166.66194095191375, 176.1485424831929, 188.37642534878526, 199.39900131899716, 216.10994753487444, 229.30355739478387, 236.1768659491449, 240.1110338600089, 246.58148622160587, 251.92069074950336, 254.926605727179, 257.2611689872017, 260.85860295686473, 263.67063242695264, 263.751447293808, 261.4462328532735, 252.073829122373, 244.92173597178754, 244.7661745151608, 245.175978261896, 245.4681907079609, 245.76823912841022, 245.83252904401786, 245.81116453385826, NaN, NaN, 22.550424072702405, 22.43679996994148, 22.95026222658445, 23.68150034651626, 25.118161992463854, 26.220981858762066, 27.246985313678966, 29.303908075524337, 31.214555209966797, 31.94263327151875, 33.19131321291338, 35.24890743453061, 35.64924562099105, 37.079411126011216, 39.502537964025045, 41.70435996187182, 45.85746938687624, 48.86923568056541, 50.73712767427545, 52.27508313356796, 55.652352577285704, 58.95738693303384, 60.348195889638845, 62.84289260733878, 64.51915234263781, 67.74580932590634, 71.12130566226291, 73.46836066472929, 75.4483769122729, 76.76283110523624, 79.11173039446021, 80.06197682977623, 78.95114833842493, 78.13610699991564, 77.98063727555422, 78.49060286295756, 79.29646536028375, 80.9896015607571, 85.03074819520863, 90.91760387744499, 94.58834449757967, 96.78632992974158, 100.74663655196419, 105.59934528777288, 105.89790397954341, 108.83293201695545, 112.51638767209234, 112.8123792560725, 112.96081395549862, 119.14037652001899, 122.10610277160154, 124.93110972939564, 133.353869011792, 142.6903623277605, 154.14935050706245, 168.51725947479483, 179.6426309798239, 192.02913275304783, 209.94339358313198, 224.12131982034117, 231.1834136598363, 236.5803572034191, 242.70249596873268, 248.28633841276962, 252.25847019719077, 256.97845853834593, 261.8572606424754, 262.7237805411611, 259.4294266970564, 248.47399714779627, 244.94113254261916, 244.9019541719363, 245.313927022956, 245.71841084072653, 246.0132172299176, 246.19993262166443, 246.1603244729817, 246.2295915523842, 246.31139158469978, NaN, NaN, 20.443368565113754, 20.183082661553186, 21.064793144870645, 22.462565079631215, 23.342817447848233, 24.44295516744257, 25.875063896459757, 26.533403554562526, 27.96383887669454, 31.198551917770796, 33.84616508306215, 34.87587870330057, 36.23286770884793, 37.26015092481774, 39.31639889910355, 42.292595423547, 45.08121069797271, 49.010161028741805, 51.800156750164156, 53.55652377091916, 55.31345172784426, 56.705604121881244, 57.50498707650257, 58.895591808710165, 62.34197085142047, 66.96524259122496, 70.11707862531537, 71.57962148917107, 73.99607432632698, 76.04814977862144, 79.26616987580853, 78.31196747733728, 78.23335453912625, 80.57436533344553, 83.13004903781639, 85.98478632438594, 89.06891040224406, 91.0530529903947, 96.63002130213653, 102.72230365143402, 103.56660959122897, 106.94582296192695, 109.305507279768, 111.65488553843939, 116.22118143216827, 121.09958591385953, 125.9839177582146, 134.1373362796916, 144.98033048835492, 159.38123789228436, 176.88896494275738, 192.25581056239906, 209.0137430639943, 224.17060859748324, 234.26589689161415, 240.11145900049564, 246.85695977257498, 253.73832415779412, 258.72758318118395, 261.1745076916491, 263.14649296324245, 261.96524130796365, 253.10829748548545, 245.46667498193997, 245.20070594363227, 245.4992328363386, 245.6907866769838, 245.89469859186454, 245.86243291492937, 246.1561133418752, 246.21839501379992, NaN, NaN, 22.734819885851092, 23.1013720241247, 23.170603221851938, 23.459058585034068, 24.33724102227885, 25.43627204997937, 26.903111241484773, 28.81104575810614, 29.91274824306114, 31.45345863511316, 33.727766652511875, 34.23391044374235, 35.11040021649265, 35.25174569525529, 35.97962997841224, 38.18064937714957, 39.86750767805567, 41.8502872662779, 45.08443595258848, 50.154292884147715, 54.26281990050066, 56.7534679192701, 58.292930227860666, 58.58110619085869, 60.99588738640347, 62.166599179799285, 60.844089824692254, 63.188570763343506, 68.68904203037901, 76.5446074798487, 80.36275863618664, 79.55499233813453, 79.69693043159491, 81.46163696337427, 81.8950328841543, 84.24048820629511, 89.08568979689306, 92.24301609340748, 98.78432879611948, 102.75469712900781, 105.64207653267366, 108.44161544882856, 111.69190697704133, 117.29205978740279, 122.46545630038615, 127.21826566648751, 133.4342512870735, 144.11034992880326, 156.1394845062255, 170.22882757085586, 185.15230200612086, 200.2435362509533, 215.98521622740537, 227.45143549633016, 233.6537589928741, 240.19540447598763, 243.9416853276101, 247.95578139356857, 251.57329600941975, 255.08781867893433, 258.28634647248833, 260.1896063677469, 262.5573284371184, 262.7571783364257, 259.0175240350317, 247.03862905556988, 245.31768453437377, 245.39154656101246, 245.686173906598, 245.98260142656653, 246.17440727657203, 246.2629822907944, 246.09739289887725, 246.1661504610076, NaN, NaN, 22.329687539246382, 22.91682014025894, 23.281008158936842, 23.79203460677967, 24.671388277388683, 25.920344490757365, 28.421202352590416, 30.408563149551327, 32.17004144515274, 33.783706057550276, 35.101678967439575, 36.64069799066075, 37.811191227911124, 38.83677290956551, 39.932600225918506, 40.88090466187905, 44.69738980636637, 49.83822949059104, 51.449924329830864, 53.06236717080818, 55.37196173588822, 58.014308245038514, 59.11192693389882, 59.88385251076827, 61.08745515694958, 63.28648030027919, 66.58878242093415, 71.09881212353588, 76.16320795410577, 75.83606968199643, 75.71795843093287, 78.57674166314227, 80.77273839844139, 82.3141411236969, 83.18922397949395, 85.49361189368027, 89.13577251297289, 92.88758870669722, 102.69687140545138, 106.02012250937682, 109.51941495285944, 110.41892352923661, 114.11712939873358, 117.97006376360217, 120.6159535055664, 128.4497315301206, 135.54355412942448, 144.41065406769843, 157.32707559319627, 174.26889795860555, 189.17194880889033, 199.61578095217584, 211.32218831218074, 218.77481768978026, 224.84456173711277, 231.32837522356328, 238.1496020255916, 243.5994573199973, 247.61261097024132, 252.92565331055263, 256.6179777858558, 261.42853786137147, 263.40804150500173, 263.2239280007433, 259.5050107623349, 248.25764755782788, 245.2544291175562, 245.44252911808286, 245.7394384177493, 246.03472389444332, 245.9961743880764, 246.0635927220529, 246.14711054076474, NaN, NaN, 20.594216389209397, 20.48273538153845, 22.176362294529586, 23.869787851162453, 24.5671932798024, 25.63137166984146, 27.286738744523934, 29.343891005772186, 31.219202370962815, 33.24226664602528, 34.1956465633798, 35.51383786142311, 38.27177888126511, 40.10768014698977, 41.17022882397001, 42.41319527194641, 45.606723854272296, 49.42769633779374, 51.70509634206126, 54.680218725040774, 56.992898363178924, 58.45656425628917, 56.54086199092684, 56.3085564920998, 57.916616857119294, 60.55667503618807, 68.56049936378884, 74.95013252571376, 76.49528288975415, 75.82715522022163, 76.85154662460536, 78.24357397950851, 79.19406010972882, 80.94755905421374, 85.05208555703544, 91.51263694119866, 95.92924445432946, 96.07801359819065, 96.24488194605527, 101.02428922291506, 105.87927171091306, 109.7438495111729, 110.97388484288238, 112.19946417925902, 117.50347005248541, 124.80136706094726, 130.01320634319438, 134.88432820895545, 145.53693474798334, 157.54512997373965, 171.45558277048576, 184.29762834649426, 195.70306596743814, 206.61319000588944, 217.1842873340936, 226.47744925031733, 235.12323892025833, 242.336408416992, 248.96657745664592, 255.3223071925446, 259.05796664662466, 261.17633100481527, 262.3008092970404, 261.7116602800419, 254.31952008041134, 246.61842703292615, 245.41261945156973, 245.73388940234886, 245.98285283021582, 246.1603229203176, 246.33371678989843, 246.35498983256903, 246.53073159873637, NaN, NaN, 23.95606631404023, 23.989673477638355, 24.35346156037332, 24.86366097434997, 25.63201275450333, 26.512279083634795, 27.429720604379657, 28.602942605035658, 30.659631276301496, 31.941004240187624, 32.30814653038908, 32.597840676610666, 33.84251269337665, 35.45732325623389, 37.18243650558438, 38.905271609817916, 40.406952123170186, 41.50385897635157, 43.52076634292748, 45.3552454056151, 48.254731930858924, 51.77819497857679, 56.774496725336824, 59.93247021895043, 60.51962462268073, 60.36337094830774, 61.45412494613674, 63.0617392551827, 64.08547851650259, 65.76955014403123, 67.82130554437627, 72.07964752436023, 74.79256062141118, 76.25463909319394, 79.70564948354762, 81.76163612990513, 86.01338731458387, 90.33712874649876, 94.3063473743711, 96.64572815537399, 99.56189548974893, 101.63705209479627, 103.99045204015725, 108.27083969454094, 112.54196535720853, 113.15291643315902, 115.37638323322832, 120.09700422735138, 127.47412747379954, 132.66496565869056, 137.0963094448882, 145.98062063804875, 161.24487716814966, 171.92349288118857, 182.19645694768022, 193.54957555478106, 207.38967768271993, 219.68431680834965, 229.21078283166756, 238.48888134008095, 244.60885174695812, 250.6423660019232, 255.62976049584725, 257.95696592113535, 262.8172346218616, 257.4096421431016, 251.1754483686388, 246.60622221306437, 245.5513375562619, 245.72607561898442, 245.97435767001718, 246.07999834531185, 246.32762466537687, 246.4295329570358, 246.5246276458186, 246.618996677814, 246.73611078352698, NaN, NaN, 22.701179934455567, 22.661925687203336, 22.842379059687154, 23.317951503563343, 24.675704763066907, 26.033449618052945, 27.281654519147217, 28.56571194079208, 29.813870695413264, 31.172031159934676, 33.70662533595874, 35.50345389089477, 36.93265782167312, 38.25270458553758, 40.417842343775575, 41.44162936798775, 42.54100366043376, 43.638361559172466, 46.75536982913428, 48.5867127753668, 51.23055656633415, 55.0466573460966, 58.57487391368802, 62.39321169089889, 63.861840250841254, 66.12749298900496, 67.2170319921703, 67.13529418657677, 68.01015308829722, 69.61856491893374, 72.3346813668088, 75.19710264647262, 76.15004115714525, 78.05690831744651, 80.91751628385204, 84.44631075893085, 88.91751325018622, 94.64793340592612, 96.63492199900233, 97.21420539845634, 96.9613870869974, 99.89266666609034, 103.58816918434141, 108.45926759255248, 112.74561469951821, 116.42804151580695, 116.87899133034658, 122.64807956263388, 132.11388364190086, 141.43729125779222, 152.8267664244059, 168.10860772102808, 183.9099399781999, 195.50048520188426, 204.66630985426073, 217.73757047588487, 227.36517878990583, 235.39395346305673, 241.3635602331568, 246.85886789426934, 251.5188871161854, 259.41808116042245, 263.38284175112926, 260.5052310187805, 254.06207998432822, 249.58707403454048, 245.5353571032518, 245.4114341026808, 245.81016946447699, 245.9108043777322, 246.2367830202864, 246.26495280960924, 246.37223612899828, 246.40927252097703, NaN, NaN, 23.775560791329653, 23.47752477766867, 23.842895291498106, 25.164278663052432, 26.92781171021531, 28.47091132824004, 29.86599058647565, 30.744668364395505, 32.06536276799343, 33.898959093623, 35.511968658259946, 37.346790849606464, 40.06533659397569, 41.822659790656736, 42.69548599209085, 43.42582651643703, 43.93593753553885, 46.13833096849493, 48.487290943868345, 53.77421648915644, 57.66545493045483, 59.93384776407594, 60.36821682598346, 63.85385543177672, 66.49688684746835, 68.40608342201327, 70.34618752451871, 72.02895272379709, 74.96119524482312, 77.7478523937796, 81.23378765932947, 83.39174221101943, 85.44750879975348, 88.16497643453711, 91.20318801582673, 94.20660556490577, 96.30255294887051, 95.28102630308369, 98.22575598946715, 102.77354085794404, 105.11457099949537, 106.61155328501577, 109.56472635237186, 111.94896371675699, 116.07275308638722, 122.57871013152443, 131.734710405119, 142.24210227609595, 156.29689355477265, 167.54980006021822, 181.7184818530178, 194.08355872267256, 202.2804380797702, 210.54781095624892, 219.85906831199603, 229.81594713651089, 236.06373298855382, 241.94263251268555, 248.5374653961051, 254.2978158586731, 259.4985977572654, 264.1872797065232, 265.9217123924433, 266.12949947662065, 257.9113825300345, 249.8011836926862, 245.48875703949463, 245.44392911991628, 245.6988636356709, 245.87473368854447, 246.05657502386583, 246.01603235080003, 246.0502915454433, 246.02146833951525, NaN, NaN, 22.702158884796113, 22.552338254874815, 23.249194053048946, 23.944994375180997, 24.161922905972467, 25.371182049804386, 27.76034885613607, 29.303007089746963, 30.329794093194142, 30.69213274991255, 31.312173653998485, 33.55034028034139, 35.535499184019024, 37.259857561161255, 39.68224351530044, 41.95730269339393, 43.71552185175354, 45.51739504114442, 45.40768615059738, 47.018605951052535, 50.767153805843954, 54.14382189789912, 56.42005475497809, 59.429465189925196, 60.15886176189271, 62.1400525939159, 64.4851745230418, 65.94606051170692, 68.81099500870391, 73.21187005755851, 75.11950617561682, 77.24803693735383, 79.81169663005734, 82.8177897021051, 84.87222603941092, 86.9962667644694, 89.76935301123373, 95.4923029132621, 98.43593429821439, 102.39843333675535, 103.27326521568453, 103.72669483748864, 106.81339572961564, 112.41810948642953, 110.53521759361938, 113.06614419005552, 116.47438023834046, 117.37036361910475, 124.32324013827136, 134.07362087680957, 149.32404691533606, 167.7517542609777, 180.82598561790778, 187.49326465821093, 195.12965590635673, 205.61529165942957, 210.34397101280337, 218.52032854244848, 229.99877429448193, 236.5002624686721, 242.5958429115666, 249.0567591764994, 253.03115756536025, 258.5476519910508, 263.6153741531314, 266.33544023512576, 259.87597452154364, 251.3883463820111, 246.08778608986904, 245.46127926990482, 245.709736182968, 246.02911642612915, 246.19679516378432, 246.2899279057469, 246.38458278894566, 246.26666295510185, 245.95719508178752, NaN, NaN, 22.811091155300247, 22.550230763791358, 22.731072549099085, 23.20589651974531, 23.866263494485207, 25.298078116945902, 27.538805070888177, 29.85645871350916, 31.14165876281967, 32.53579369084716, 36.064336827922624, 37.68245335918822, 39.516267465580356, 41.86292783212553, 44.874409798854664, 47.666032259286766, 46.63580792350133, 46.58751304819953, 48.08888293196473, 50.65456742072573, 53.84368415238368, 58.61705746820431, 61.48057047639599, 62.656032376501635, 64.12348685306452, 66.02730417009961, 67.85410242903701, 70.71682317207359, 71.15302222073127, 72.98325982790023, 76.8677748448968, 81.12051443756317, 84.4862051143052, 89.0296772891143, 92.25196477441762, 94.73740440327362, 98.1854198838906, 100.470888462106, 103.25929320290177, 107.14453695512339, 111.5817201395002, 112.31190361063022, 113.65967680714893, 114.57727046704166, 117.39256120414191, 117.85607746351499, 119.93560419022076, 128.78827369376208, 142.0991039819568, 158.5549788420761, 176.6773439556107, 191.15082167713047, 201.17777984842434, 212.12272086778046, 221.4768695696239, 231.58043396698952, 237.62257099704584, 242.5306275285077, 247.77745999856955, 253.81198985177457, 261.1113390812844, 266.1039878872576, 257.03281054271133, 249.00381817514025, 245.2816486051806, 245.13137526884466, 245.41931327519728, 245.7158997767384, 246.00684273982546, 246.18437964723356, 246.25393400347258, 246.3141319740528, 246.27815348608218, 246.594541137162, NaN, NaN, 22.221808082236038, 22.329438884222803, 23.025482170629775, 23.75804081699179, 24.122746647504798, 25.002701681751823, 27.317611610142855, 29.520778111567676, 30.80414799976653, 31.68355731979603, 32.631993302315095, 34.39354660090651, 36.29826554911971, 38.279244742620186, 41.06622407685808, 44.51515574976891, 48.51582574959973, 50.162271033359026, 50.529207889975346, 49.6768835003911, 52.75963778499417, 57.825464153879715, 61.639877690005285, 64.42727682949428, 65.52490265788774, 65.59275749066974, 67.57023893207834, 69.32645071876794, 70.27626165182814, 73.27865482458193, 77.67366475874209, 82.36808478421811, 89.8585601696564, 93.75802384474935, 99.1899503192961, 107.35293047191335, 111.8393797048311, 116.04811234203544, 112.16717543198547, 112.0037984671173, 117.69893011512899, 126.2474030864142, 139.05297977801, 134.1110369331247, 131.18002704207393, 141.50273357168118, 150.2566124548507, 164.59795022449293, 177.92115608398527, 189.30859156391426, 199.73347234773158, 212.04686898371938, 221.94911452111103, 229.7523413804016, 235.66114233279856, 239.90447141022975, 247.76371069309505, 255.62697302824208, 262.4191143443135, 266.3195747279826, 263.47510949962117, 253.7732533829319, 247.34082924923536, 245.12626791288258, 245.18864945808505, 245.58959659404, 245.76570903652689, 245.94823794095853, 246.01478896254045, 246.07326924209738, 246.15377670178717, NaN, NaN, 23.591080967237914, 24.215516607006165, 24.91170823341797, 25.129495232266137, 25.309699266606923, 26.11387428572898, 28.576134283750424, 30.37542793279396, 31.844455911834395, 32.94323464671442, 34.004775541585545, 34.772435147479605, 35.65067274368298, 37.44776111632004, 40.01628628476257, 42.810371632066214, 45.15835789499984, 48.61370673570636, 49.826170291709474, 52.10377137141375, 52.870526008742516, 54.77252361544459, 56.68117034338894, 57.85185978462884, 60.935967172386796, 62.539849602727045, 65.03531351546539, 68.85023098439159, 73.40105546615895, 78.24174619444975, 85.43337590019551, 87.63928568790946, 85.8710572148636, 87.91914993282809, 90.55105093437886, 93.04682229943853, 99.79982165449785, 115.22497750793741, 120.5110951287009, 122.41607818246582, 129.5269169762119, 135.14377935238974, 143.74331533903475, 147.7237682052739, 147.41620535854176, 149.61570745753477, 152.95694265184952, 155.770664460264, 163.1276875204356, 170.269369262345, 175.1615600927909, 179.49868218931343, 183.8427764884539, 190.32841016057208, 200.1722828350844, 210.5870347847899, 218.21351261920523, 226.3799234657936, 237.16495845250407, 241.85372475002688, 245.1363709088037, 251.03763567839857, 256.7865883955169, 263.0201952889185, 266.37552646404254, 260.5679119485362, 247.9904758850942, 245.18507237575292, 245.35792317743096, 245.64428963560368, 245.8156291738461, 246.107387361752, 246.16757478522072, 246.22753452127372, 246.30135657278745, NaN, NaN, 23.183271044647274, 23.03296872563386, 23.87675569481782, 25.052576573116912, 25.380119055962982, 25.706804517815918, 27.026908494024394, 28.790926299798322, 30.260104409241524, 32.05853321064235, 33.453791000969595, 34.59071055726584, 35.43338834941922, 37.0097127647621, 39.90845230098525, 42.443065675353665, 44.38585183817713, 47.17793880487291, 49.93506075164461, 52.68552616634514, 53.963320318365376, 55.94182486638524, 57.84809194313208, 59.97215127184957, 60.69986838927468, 63.41703524956662, 67.23414049500332, 71.63693381571673, 77.9484518960289, 85.65536187973954, 88.59041072611714, 87.26503233388, 90.34877556022215, 95.26362250422171, 98.85410554495803, 101.56559372238627, 104.79113051534685, 113.08108814175138, 118.58536645234638, 124.01047812225286, 127.64111944312278, 136.17506520431215, 142.13791965432, 146.19458050658415, 149.67938808714618, 153.00663879698595, 160.20237726078958, 169.1679830464372, 177.84139014719312, 186.51449831470546, 194.17829454786246, 199.1491817125678, 207.33250044614388, 214.7179634919651, 222.96000365138488, 229.76456759227185, 239.1993226693374, 243.47645237493273, 247.39952261408598, 251.95475470889363, 254.83957973830823, 260.56594182842673, 264.7996140068545, 266.141141775596, 266.85730823324064, 263.2364620740722, 249.83030740129402, 245.14161820212215, 244.9506759291916, 245.19838897628065, 245.4513921940312, 245.55285601723594, 245.65209104328372, 245.61155778378114, NaN}
    DOXY_QC = 
      {9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9}
    CHLA_INSTRUMENT = 
      {1}
    DOXY_INSTRUMENT = 
      {1}
}
